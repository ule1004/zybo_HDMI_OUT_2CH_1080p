`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cCEySlPsI4ejBww/fqs4UnoqE9UfouZDDFSjb4N3sGLEJ6+IwjhcZIP8Iea5fE0uJjk+odCZCK7I
ZHPiobp9fw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XFJ2sA4LXRB2zsXyilB0EQfyEADyEfO/Hqzlh1Ynsjv8lPUSfy9WWl2BZTopm2iMNbGfO6kZH9Tv
xAd2BTD+Tq6NnswiY5UHtcQc1XajnMFzBSMRy7QtH7Qa2a1h/TCedr3NaFObq10Fosdl3FN8DIHM
HsCV1qNt4EQSDrCxNB8=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F85bwWlrEBEVbF5BTBb4XPSA7rP8q0rR6/cAEfrCB0DmUwjPOava14RHexa47isokAcR9h9zkGIU
OkQ9r6R1bpWU5BLZB9IkpK1iBwMOzHOWkt2T757BthMNINjl4fR/VEL1vJaWbY8xxMZzLqsmEsVq
1Bfyqi6xaQPeqq91yQc=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q6/Wye+JLvqYcyZe9UdxzhGN05ktzhwaEcBJfk0knDJ4UQ/tMCEDVhpn3e0H3sIgE8MxvR3UuqHD
LqUr4nwrIVxAh6BZSghtNko2U7p+tc2+dlR+FudAgukdSAbf6EhWoznCF/TnpwUo4bWOZjlm44SK
blAUmlyZqQiQ/TkV1BOUHsqudqXRNbrXlLwrA73iD+aBED3JMy2pO8G26zIm9cnhIFPOhnDAFFOK
OoP3vVi2BbM5hk/CVwXM3WFBLO36phGPwiAIEhc4k85P+qQO8aG75dWbjY6KYeXHY6Vk/8zR6pST
r0H19YpkySQahrw5ZrEM6IgKs+br0FvvZz0wKg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lg6W4aLpLtAJ0i5y9EjsG8olD+g68hKAQTR3fQzBg2I0JfQrFz++y2m3rKh0Som6WoxCu4iuwNmS
uu8RzHR65XeuJ/vs6KITXcrmNLtDyhGQmS2KmndufWl6soJy39giQ2GvkK+7TWt6n41tuOi3rq5D
9BrsntuuZU2c1+NIW+nbw8QkZvH8gV80SEA5FC3aAOHN92KfL9SuEYlx0KhjVDOsx9QZv0ruIWob
kadMURor0STEq3sjMZDZlcbbMzVOlsm4EqayPHDt8KB9c07qSvKUEE6qXRXO/xj13Rba/REq2O5s
jqeL9bd4i4qgqIT0kS+UxPfsK/lv7ZaEwiuYsg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fNJPh73T+FOGjOEMmwSs3zJTUNisWFXpt06qHONiDrI1LUgGG3B8wKGZuDXSoujMw5W2pceYrjuT
qKVrY0dPRP5tpEd5OZF/OtQWK6qRTtMV9Zcx0VKZSM6krkjJTL6D7kqpe4/7wbV9WtbtQ5l0Eo8d
sAobkGP2bNR5+3pRCO9xSSyRXso3vvibl6g+XTOykopmPzOtklAbRxuxwpzchG0N3VFXm7ofB0Ke
dZ94s1B+cAK8bc9dkbYK/WgUhsVJeL9N+d+OqYmHYMpqyD70Fr1vCpYkx8kt/Y5+aWrp+sj6kvdH
kYVt9NUorW965aCIs3YNxPH1iqaktw3mMyvs+g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 270832)
`protect data_block
7wK30RTHliBW0nhFOGMAKnoh6UyPx8E2ksbVsJM1NEGkq8nmY+A0L7jWqI6CCvTTmxEH8NTOXal2
6kCRYpXo1pFzGEwmApM6pGnMxtS/5GNPfAPBU6Ks8sJLJrKPGadCRiezsCAVSfiVhDoRJ4gzEJfR
MsmSJSSjUWXY5/ONmoC4MYeK8micech2JW1vDLn/ann0n56jRDsE6EYcXsXBKNRrZ0Hjs46z0zif
+bWWhzlzfQy297lflFxnQE1YOsAOFl/xK1s3vzxdFobNSTY27x+4MMmJ+Z4SegSgAR2JK9CH901x
cMVXMahrY8Iw8L43eVpuz1L6xB6lvu/hWOup0F7yA0NM2GRUUtvjV1ZsWchREHKwnojr/owe3gkn
Q9idSGTmBNC2BuF9kx8Ix4hMqtrzYvDfN4/YXC7PpkwN4c6IRcXAiXrEM3WBXepfWIqSTk/RetIg
G7c2GtC9IhRnkEIMcQETGKuDENmdrRUqk8TN3Yth1hzUna5aTT8LO5UIF/8R9USXMTu3LGaKXbT/
YZTsrpERO3FjgeOaxWmD1A2V3H6jPguGnys9idj42deUzqM3vnBTVda0ZB0uqBEl+eMyjMDjAsBp
xt6YqN51t3VCJI6vvG9De8j4DE7mC2K91DUPHOxMfzco3at3lsVsh9aHP3jfXVCKesshQyftXgbs
PUOUXPBqmAiGvK0KdA2bu4sWvf/E0hq/9ipBpOttjdh+Dzb+IGnXAOS0pFp4w5UMfFtP7aceEloC
7MxEjSuN4hu8W0t1raeeOZgcpZyp5pOtmUtY1g2PuimCftzK+aSHq7MbIE50rMPOsgfGm3KL9Z24
wwJw1Z/jYzuhyjJRkuaZseIaUGCn5AP0Hoe57PcHv58ZYEQvqEulZvevYrVYwqNEmjtvl61fIrdJ
leuYr+Cry8saNGG7oPWTS8mzgcND3V1+LAzbYEDhwrpcasTWOlXF462ynxKOmmVFEQ9W4x+zERS1
xyM0vgb1pFNaSVKhShFE//N2nFZlCD2dmlPgxaou0lppO/W1E015KB0hLyo8gfnfWCCtKoaVRPek
FzJOJzW2ewA77QWUtfJhDHijGW+tQJhqZNlSJIr01X2zUnytxI/6xGZ9UuswjLbqnczEIsGA3eDu
njLSbmyhdDm/5TuuyWC7v3hSotqf5vg8aAJYORWujEYOhWj2jUNxTznXHTsKPn3TbWinpFOgDH6+
ypaU1PyuhI3Sgd8biRWFx5O/Xz7E3vanDtgniOi2BiJikxU8SqLPd8I6aqmDSaXKhgHefHHSTDez
mWQStjdy0JwAc5fZAbSnfISgyPQnqVPpjEIhJ4MfM5/QVg11IuIx4rVR3PzRPMquPxzZr0mJu6v5
rTmXZzeil8AvCDW2lSRH1Ezw29k+dp/Sh2VjP2KyPgHyuueJJGFBk8a0/PPI3K9fz/pO1DkCfqpg
UPpmN7p73nOzcOGpYHcZilBD/Z0z0RnP+qQHGj5GqS/EhdwgzUs9ecRUwQOXbuF0cpDCVvo/naib
ipX3evwia8NP4zX8ZnqsorIinsXOziL25I0zB3piVfPje15Dl/h2WoZBWq57omiGatfEJ1YYJFfn
OJSMjvD57W947R41Jq4Dpq6Mps1f43iidoDv17e1XHSNHbrptLsRyiNTCrVjARr+tv0KnfX0O+ch
RQ0vk/H1YjsZgd1wG8lmrQjzRr8yv8KqBgvv4A31Zk6987YefM3DNwSzSMB80VzpeWd9Zi/VAjcV
TcCb0SH0Bt7ukY7PpjeQJMsyOCUz0Nvg60TWkZc87Ir4fY6I/dPiujFgMSi5bggRc5ZygUyZ/ZeE
/zeSGk2snknj1XYqb6HPtw9GSnU4owJEShx1Zpq+/lkMujKuPyBU9nr/9Sprk6a8HQrbG6M43lho
isqTxDAwdgfX4cy6bTwtv9j7Tq4yCylSTYiUwxk1waCvioDRHkbGIfa2teRv4OhDQeyESLycKUsS
Yl10C+1rw4YRdCrw9oxxTG2H4rwgWt0ekvE8hPymBSNhMvXA48DDdFc0qxcb+fiKRs8XPHR2u7Jf
gwb/qcoW0D3UJlMghClsm2rSiQHuEEbD8cpplsAtWKhlHHbuPt609tQOlnP7LFoBRus+/K1IvLcS
R25nsCj6ySZbccYbNXTxalqgplNdo/GQOHdMtQM/+5yt9RDKGKXGhglQikBCdP3ZHLqzbZOvr9iy
4+0sXFIdfGSXWRFoPKFuIzHorzB8N3HPgyB1hErMk9/KKcabNW/0Y3160VpjeHhsSEtg+p9hbIbz
feDky7BFJc2YDPaCq7NT2MjmLVwDnU56FixYm+ze2BGzSoTI7/fv7EINGXVw2lckuVY0pQI1K7h9
CCL4qaWuXA8HlslzuE54PB+vumoBnl2N0Zg9RzO0hFNwmJE59PYY+T7a2uHePJbIY2oEsgXqRfxS
UFj7MlKMbec2jtYWNfNElvxsuaOGQYKFhZafdxOgZpe9lnBEPtG64N72J+dvFT3K0xqRxQMGG+/l
MHR52apN4nxdTnTvVsKaW76dZozqyqqTJy8lSVSX1UfrcjyLLPHNkHyE1JR+oYLH0Txxac0UtfkH
ylhzORBNHP3ZFNRw0k1BqiT4XZCZ616tWQaGocLNpi7zfaH1h+StoS2rUkr3JPmt6tWZDnz1FQ1B
ljBCNJsF5M/TtYWnvZQx0FmM7hup3sR+EI4XZPUqu5TwismHhd+N77N3XXyLOdKqhLJi9gK19pC6
rFQQGFr/P2YvcVdCseaKdiodRr4FJzKqoD8KeB9dEPv7UBaCOeq60XzbljmlNaxAhLqjFnUOs4BW
S5Ri4DMEWmHD4JKLnGxNHBw6uX17DVcsIbTUQ9YJI2mRmEcJC5tovhXwzMdjjVaEt1FiKLACGyTV
4zvpPpw6YFQ0WaEaQ4V/OmbKjBWPjYhPDN4syOAG/JnEIODQeu+qBdPpT2uqkJvig1DncaUlHn2S
xxmMj3UmCgAwgqV5dfLGxl/vfGN6CxnA9+EAwQTjYvv8lvq3CfYpQUzb7DTvPCrjexEV/vf9Ady3
NsP0vreRnymv7qGnc6rQV7F3G9RwtXsFUFDg0K2m+s1W82BzdCIsmakNBwbAgh6yyS/LbyqgEvtZ
YX2i8eL8+6/s8/h1vedk+YaX4JC4I/3TO1oPmdrMPvFJF0PSHKb/wXUtVeWo8567H5ReZFCt7B71
LKdLUf9jxYVAwixENvMKL7N1JwprENQHmxs5+4lWaKkOsZYxbZOHXJ3mcwX9hGlxi26ttg6V4LwH
s8QUxxHR5KSKuffK+mhFyzHg8IjCy3gcuEhWJ4io0gUMZm5WWmDiRAePyB7ijdRT87S3qTPB2Sgi
isV/E3X3WxjrLwlwo14fuMoy8jX7KmNxHJ0uHTsniXYn4b7t0TDNLUy9i2fuGow0HtvsE+DeUhGm
Qhg0E0uzl1wHcsYJ3Ze/6jTf6F1Ix3IjDki30iMd6qkytDx43pToY0CfPS8IkS/fQWpijpEeHWnR
4xG0fTVw543QG3zP7Od27xce3O5rICYM6+EyeKssGFTEecnc3mY2dv37SAuPS6Mtf7Y9to8M37Nh
rL/G+rI6IRMYl/lg6p3geSSLeqraQrJHhUPmeiHLfFshpyFAWdlJETiaw/hAZgPrf/Jl7XNuhlLX
saspX3/zQf07k4krMjB+pxeuyCF1Bey4k18M6dJ5mz7HJVs657YlizQjmXxMYYKkH7GgtFijpg8b
Gxcsz+Q3km6Fd0GcM8d9Nw6TQ5K4xVHnkEh+R/MZtyklUnHIsdYB9ORzpQggWsgxHcSluORDTCwP
j9SQ3OmXSENT3TA1CrAhyO9X+A78NCdkdmivVYN6f0z828oofqbd45vv5pQyP2e8YJTV2FLPdoYV
rRkwmyUYQIJEnuV2i/drI58wQHMQQd2VIUW2TwHpRQaRPGmU4ulTXu7OJi3tGYsii7sGtz05M/g7
fCRkubcCv/qVaIiRBxj5NlL7g2kLOyPIZTImip6VLWjq3+fZBplE5BZYzVZ0E/594qt+Pip7biAK
3BUpLg1InWJ82YRKtBJszIhNaHr6rzOQHl07JxzKxDr7s3fFa9lRn+cPMAUHpQCheXZJJPgBd/qj
DrhX/7/4JCDKOtdZAB6HETvrIkMPz1rypPuHq/iz9Wdif4MFvP4Rff9RCK7qFxlYibIHXl/hoR1r
vqvYPLC+bmb6R2FlL3ZjYPslKr6BgEvEYw/3/k8lS150qw1ydv32BcC1g1t/8ftwocVmshf5aCvL
ocHfTzbcRxBr+N6kRFkCEah1nJ2U3iY7rW+y/LTGletRsuZP5VJUoPhCcp5l/An+zL3RfP+AajaO
nBila9+HhLu+ohfRxEzNZp7jfmfQTNxsJF/wskAMe4ctnBxPLdU0lUNCf2rlpiOIbc8VMyq7Xmz4
LmrFse5ND4RzuvD/JP5gleXdV+HBK/RJLk3xMcFiwIcMA4Nfuvct4EiKcxG3fYnjKXgP9+BXqhwU
XfxNJYR1Li27Rv0T+9W8ajLkTmSOZ7nT+cscxfW8Rt0HbWY1eV7Lv6YiuxaPncrVr/rJhRQkaKw5
d3ncGs9q9eO5vBHTBMezA1kPj2DIPR/8OLeo1E1flZUcN6z2gtILReLRSiIPY3QuwZIadnahcpSK
lWrWTKCRzuLJAXpU6dos3qltND27DTN1Abef7d465q0gx6TBha3MEYaXt4rw4j4d8SubVEdMZ3Qq
/wdmx+GgZy/1w3bG39gv9ZBM6f4eIyYYTH1H5shfYNpjTFjNRcvoeegBg/U/1dJHGdd24ydxiLTX
E8oKqAncQ8prgoWgiwA1PK2mEa0tYfKtNc0MU29D2hmcpcrSpDcPO+r674v6paGYiwqRizmuO1vw
LYBwYdVnJcn/ayI7X4RdajmoAZpr/jypZyxH8GUH6T693Oe4X8EH0qH+30hVzbOqGTACquqhfW1v
DJTo8GSMnVVba/xdT6u0DXh1yTy6wJxtI4MLZCuCZt3awCnZdGU63xVufI9g4Qg3GM48m/+/OWEM
IyDOhyQeBnfO6X/SJLxcyqUziOjScPgZ6FTxv6Efv25GAnkgSub08L6VEF8eBoeppvsSFW48l0S3
yyh5lARXSS66tiwsoOrgxQHMcguKEdG/fsPwcRZ64qTWrmQN0iVuI/6KRPOkPl5S6cbkvV/26rD8
jqcBFCejxAHx8r/wJ54Nzl7GraKpMQzYpLmXS+I/npskhymNj1hAZ9MZzz7f9yVN4JoFqbNxT3ZD
6bOYsJ6T0seXht0xwGotUyn56k9sIIyyEHXVghFB+9j4XnfSjtGRSvl51c9zeNaTxkpffSM45/ao
nl35aCPEKE6z3Fk2boaOQw67StmKigQ/lYzH1quB+4tpriZo9jKA3Wwd/XjBFb287wW0uk29qE5/
lKKCtczVrUBX9Ib2pfjHAnnAeiBlql9QJBLwg9sVsa8mOdB/7VwxFdyvyGnw+SRRmSYIZBzfePaD
AHPAcwt6Lp+coDSxbcMCNYra5ndm14sdLy7HwLXFeYnvWIa27cZQhiTI2T1yrZy2L+m2gb8tzj59
QY9bzeVJqEEheLiGVEgbFPac3R98o7R1Fwexcc4F6ZCUCI1xMCsmskX/DVCDh/mx/hOiYdYfxu2T
YxLIBHBdOkZrA0Mcfd4CpHHk2gT4gQuKy2wqN19yot+h06ha+7Z2cUr4LqC0toTexCTAM9aShf/a
3KogeIExNEs5WgY/IfPaE16CRwcLyvME86KsMShL4iUE+CJWi7ifgFu2q5CONALjcz3P2xXr8nS3
tKRrLU3Fi3OHwTfuT57aIxRxldfb8QwGPm/E0JQEp3evZOC11iRf28EJ83EaXlmgDPPK5ph9q1yi
4jIyenPokAP+XF3P/J6+9OBCmQPyD078HppCkpcXDSbrUVxq/Gwprmm5l4i2DBbJNmvng4CX4Q1+
eCgFheC/kbGr307YWDRJz3hDz0/cI0smULLiuis/r5eCwLwoj30l87cne7PXTVyBgLy6Wczd5lBo
vJs1xNo0f2DS1L2BalwAOMXZ+n6nI58MEdzVRjMJbWhOyWtSD8FkAmrtLTPA9W759/qkI/hUqjrv
aWqFFTmXt24wJrD/B0jeeC0+9MyclCfFwDn+hT+FtOQHG9zZOcEt8ZochomiG3wvfDP9lr7yCj70
vfCbUKWgBKS+Dt4iloUKnqtH4kzZi12YicPFGy39z+tEMb4Je0KbYTpbtiOfLG4AIzh3xLz0Z1JH
b4YHc4r2DpRnLdhA3dnDWcdyUo1SKEg/PRY9aLaoUl8DHfGxcCyCnAY5JOnb9/uFVQZKjEQlBo+n
xmuk0VWEZBzBsJiJHEqNnmCCKH4uhb0UhRzZL+kr04wGm+wHxFJUx1fmH1pPArdN/LMCmiD50RDx
RhKgnZYQ2UvaK+vYKtrentRkH42NUcPipMAx/MNPsoLT2BkjQDEYeVMOqqS0/DUHCDKtqnRsyMPv
3Md5+ioFmV/tbIgWmUFDgb3r1T7b38dJTf6Dvy57XR7hJPZfH7P07abOLo8fiqMth6R3TZKT/1Rd
Ksn+0WYzFLWUQisOE+rcw4aYDkiRMYbncyWZ6ZgvUJNEAd7ReKVBhBzYtKSyeDUEy8NopD6maepW
S5h1FgHnPo39Kq+x940yPVvtlCL5OKneCOzmhkfpBQJoQzlZuR9DGl0GRP8xVX8olfH75sm2Pbnt
T5r/fFEygNAT8OP4wD1U0dTiXYsiGMJwloh/CPVX2nwQFUOMsvCgfSwJWxclbp3XKsyjxIp6USr3
0AHm5j1b3g0v0VphuWHR4Yz/dsBQ9nEMsKvAel+yoOogmi5TOs/qqv+8VDZq2y7LBUie+s411oqX
YMv07v1ZGhl7uLKq/LX4NcEOer4d/QlleF66ouKbrR+hRD0glHk9CJYlfuvW/RUa4jTWqsp4PGcg
tPpJhwZk3XvI8JmF+aq9pExiKF+HQn6vugKKhJFvce/Z2H48phz0TrhRs3ZCI8ABJbnAWGp9/JYo
r1KmZI38tvPGTw31K6nz7E1P6tjX/LIKhdzH+FH5v4sEVY8q4O7aSIb1zL9Ja3YFdTTjeYVhVk0U
aRpzoTwFCt8GSnPbL1UVySL9OkqCe0AZNpykQd+Tr639GEaVI4MAQagGogg0BcGX/gpBJh7uR4H2
SfMJ0rz4Wtt9Mwnja8j9JttjVLN+tAWQZBOHY6b40hKaoG0ZUObZbx5g9+q1VRLb0tIWLLTgdL88
zlPk/C2YfXlabXMI90wZ0tLw2OuPP0YtmuR2aD/e4raLRwWJ3aq0fPGaqXAXc9U9qg1IWoU1EJFO
itQ24kcwe9ZuwXalpUmQ0w6cXEqsDzXZpf3KgiEYdfnnRue4B/T6w0NE60i/m6whd0yNB7bLnLPo
xBMAhff0+Q/DJg5+U40f8061IjkyPo2V9tb7s8nm8bBmcYWk3xkUlr9sPE7Mvqh6LyMjKEd9rBRz
FHMDqhgskBYHxLoj4lYYpdKGpjNI6UcJ+cVfuIJykMP6lzRrzQmqcFG/0k9HlVglehWWjzrnb5qB
A32C+GAOV0mTEUmc7k9OzqK/XFbzzCLMVj77ejb6ab1knq13XyfX+bPf/nJoUi47AQ7wkL8NlMgN
Y44U4PHmGyoZP7nazepr3AeAjUW5IgSu+oDFiuHrNDAbnbY/l6J30QcOtDjOP8Xam4of3/7zkD6V
GV9dW5/gUbCm0dyJYr2Z0mQQGpa3/Kv9ThGLiyUG5j9WaBG38FxW846NzQI3THzS3ActFkV5u35I
So91xHPxD5nBdI/sXJNNAWLF4p1kjm1oF35vTZTuGLiXCoZIGQa3Q8Oabsq+b0T4zPMCIzn876PZ
0qnkxDaqEc60mEaTO6ox0c1QkBiKEcvF2QghluRXc+fskSP45WuQ/LSE8ZaZ/pMb4EeZFCWPNkej
Cz797H8W+8/m/3n58tqn0yC1KAiwaaEGg6oSXmnDG6GoV8NZmafQJ73fKOUeaO3d1q30ZrZXP37C
Ioc8D6G9mgByNZyCdqZShCtdRCAVZcIbYElkD3Fiq0JmIgFNDT0vlH+Pcdzuz/CZvEuIKObK/yfR
Ryn0yuiuTphcDDnhrnhawk0o8TtJdpWnyHOKdJCsnuAj6rBx2Bu7O2KWhwjlM7kf5MPEwqeOPUIb
xfCxaC0dmc9IJwa+Xm/MCPCcGQid6SsOCjk5+36IbpnMignagdKqa+CcSaVQQ3+7LaQ8tHB3CRXH
KK+N9ue8/m3CC7lf9bk22XoBgREOCoOzCTILGlsQgIwXBMVXqnnEs7q80aRVWXjM5hstRc9i3KkB
g1c/ZABPxSzks1kwSvmMZtdY3nxySIJ987hwxL/hJG+kiIbhPXLFIxJBfC0Mw6h4R24dSsVhsA0s
79sV7AJ90uyJK9Swe/ExwXLntX/dE/0BBw+NExXq47zegBFbbyg+1S32Qg1ziMQ5VT5KbNBQ4vrI
sBMuO0r8OYT57+2rwK39yxpnQoqCH16n/pq8SCKCLyAXQHi8Xe6ncqs65GaCW7NO+X/0JxaBuuL2
SmNxJwOU3pLtVuq6pAzMNYaL5ElE5fyWkpfDWtHb5uubxtChTY+XfXuIIETL9ayhAj3dGA85QnEY
PCEFEuxYkZNGijYI1+9EBjdyfrBzhTFRIJxgRVzEFg5z2y81uhMXNkjpSG8g6fvNFp8zaVL+AQ8S
Q0VzC5pubzSGliIIcz4W0XDVZDZt3AyYHl9jcxNS2262FP0v+lehTvsfjUg/yZkPC/gxlO2VRgfG
4wpEsD26plA96Te/ZoyiKp1dFQfkemlU1XwEhV0ZtSVeg3c7uq2UyF/vcIC2GBScjNuvxukQspKv
5MdZqQn/jbWf+VuONjFmfqJ4oAa0ayFnSBaKgHyukcBUnBv/rllwSdrdTOILplrIouDyDpgWilch
dUpf/C7Nbme79c+5FBd2GOAoFIQJuzZCN1uAyMR9zTnN7NyZvlFKbnVusrlY06LWUDxEtqmOv3Bt
8WSviLSByEnVycP3ozd+5L21Ntu+7JYOa8c6edN4hsSY87P2LQ/W4bYw3hX3TIHuWrUTRYxsNXnr
c94dkl/IyFUuvpFF4TPpQum03H8qArVu44eIh93fN2P8fY0pip13X3x2xDY2SQRir8umM7e8RLz9
lfODhGR5OaILGzzxpEYBqc4y6NE0QPx/NWO7+p/F3enJUjg/AiL4ApsBBGLXe6gOmT2/KF25CrgO
9qqIIfzFFOTNL8hbHYJScMo9eJKeWl2Vv3u3dNbWRotdX666EV9MPf6Dv3GIop+dKt+XEy7fqdhK
C0uy0DaFlotBz3pmQvekS3ZHOlb+azFKHJ7CjRhRZ3ayHuqN3mvPtOsriYwROp4XggZgR/mYooEe
P4naxSsSavSGtwd3pZsz8nLdUizlMBGte18PCZUA9e+Sh/0AvFd2CyWjDlK1lx6jszEhJ60ZlSf/
JHttxpG1JTVo3P/mJRc+bZfaLiYpTrzeAdaqV7YD/xCKLvswwYXIkI3o36TS1O+1i9AXBp87VxRl
nw7OEZo5THe14Ajs0Oa7AaREXPkwZgkqkJ3XQJZRFyCnZTPUYEo52HtmdomQBe92/Jrm2zxxxTBo
dsDjKiswjISp9GlicIJ7xoHg1hVO8oS5OE/uCr8+5fljGwTRUE3yZPro6eqAutCvOfeLmODNI0hi
dvZpOm+EsU+F/5+7P5naJ+TL97+tnypa49WR5ixsnG6+zbaV9y1R0d6fa6aPkzOXhLpg5bvN/MqB
9rjZNXDAgC9kFVKEP9Eh4ZnAWEgXHOlJMsqtOecoedWNU2KfwvzFM1C9u0o2hb3JYqEYndiz/9BY
6BVFj8fa7fTF6d6jEPaDyp+AE/vMs3wysqIIUkvyUlWvWgX51bJ/O9LrsCoFjADwOKsO0YcAcsec
EiKWpnA3AWqIzZMDwxLYNCmFk+VZyOtxbcNl721YBkE2LOc6VPVMJHPUxqg/UO9j66FBprm8BSDC
0A0ziDnuY4ZEC1C6VAyJkAbQB+HpDBCcsCg0LJt2UqoPgLFXfMXCNErUXRNZCa2QLRoBrNCrAbxq
GPDTJJDLhEeqlpUn0hjBToRqqR/zX3Z5BpbdVlD70o5E/GO/da3hgY5pdSUVOxBnlOkIFtQaF+yb
MC1neqcnIvdK87Sx5VcJJOt0hCq3f6OoR6yIfEuoWesJI2Y2ZcIXprwvBaOCbjaNM8y/vmSnAWLK
7cEMy29GUrQPhOmp+2346+iIX/OUYmC6IQWOPlN1bSmm8RILv5kr29r08M5ULpj4ODPmGqvCQxOC
rNV8fO5pyW8O/Vpfa3KyUF5ZRtNh90ZLtyf90Q/9gGnOmF30/riCwJQIcC6F7ahPFQoLKVOntrgj
OdBhOzn58b2nDdWmHywFKiwjHxah/NxEYkxVczwUt9cUYrZ6izTsU87hZJBJSJZJWcOiE9DGdYzi
fo+zctq1DPi441wJbh9HR0y5+p/4HTawqlBO7QldV7Q/FuGCeO9mwxGTpsFFDlGkstK+BvfJrqjK
3fSDbG8B9pS9KKytm9gqClC9XAIrGHQgn0VTp7hhTEptiLeLu6cridCObmzv6Hj4pVsqhXBjanFD
XJtaNKL26BIe8+6I9yZVKrvTjsnpPusH3cF65baf7jv4VyG3zYzp/efLphFUqXwfArbbDY7n/xqX
FeHYVE0OefBXwRMdYKoftpvHhJcAM5SRd+kJF9v662SPiksl7stkdgV9tmVEDa+hcYnHl9Gq0iVQ
chhcL6iKs9l0uAtjbXzQEG8LdeAW9rWA04HYSWSTJHqDqW0RFy/oaGm8olWh+3Ly+xyjiOPC0z1u
V2deICUylKWQUmsbIX2Lo1Yxk30Ynm0fo55MsBIWkBBtoF27FAeXKi3Qyn1tfyawPKw9fCOOqWnQ
OlN5Yhp0VppTtui1OOGjkz2ZI7esmYgE0hUQYddIKghiUaVMC1O4op4821jpQQpJWXrBp1HQICsx
5v8RtIdSWIN6jWvBbabVp3YRK0Tw92S4cqTQcuMsQ7mrCK9ic5AR+R59Y83te/wgF2qQ1r7uzPTM
TMoWjdQ9NMnb02FC8pPGmw+qN8SrLpw9ofMHo6+4KzDU7QHS9EDVziMoJgQgS+p3HVtWa7BOl8R3
aw47arlf/tX5L3Pwtk8QSuACZcdq0AMnTV3Sx3vZPMSS/U0cuA3gBJrFYzHwY1j0DpuzhojrFE0v
aL8qvfQ7rraC7NgnFQBAnMGEowrvMT99GsJi5ykf8IRNEh+r6JljWmr6Jz2oCVVUwMwi9X6QV7Jb
grpW6mRAOqruBVdhzm2DcRkg8SFEdnYe/jZoVOhAwhLc6FlOXfv0OS4Wng9sTid7ncVSeBj7ynW1
P8Z5AtlSOx7m1U6NVMGVBOPAUv6IaQZp4wgo4iNfdPvI3jxtFffRQq+s2AwLqoO+V6va9HsN4zUy
AhVqXwLkMaQA3Nu5NQwlwrxSw2wu0W4xxSJXq2Kjf3sEccHTUWtxek1bETOZlvPkezh4a2bEGnbs
D5/XJN6ljXugBrLTo/lniyAdLjYw3ZXATo6TDeD/CY50rfTRl+immTn0OzYvlUpaUYTk9GgQwnb/
v4sYRML82mAT2gJ4vtr5s2VFR5DV1Iv1GB197gCMMoyPogVsn16l1lY2FtTw1i9wQaDP1i4ZZq4Y
jbOrW2s5gA4mMV9bMl3UjJJO+/pHuzyZz7K3A1Dg2egqfvLMmHjDvcduzLuiyuH81m/Xp2qneNOZ
Fdiy6FgSsON6iJaV9mE7bhEZ1jAOkw61UylINLNimZQ1HDALGHpK9bFXhRMG2SpCEl+UsQwx81ja
4BnATydl81YxZ8fZBeIH63zrYqqurMgJwJZq7F4Zc59XxdGG6NUhOIcNcnDH1pzhO9w7UEVNDmrG
9GJmLsrxcWjxyariUtZeB6d3K8bjyIucdQieP0+dml6MGmgfUUHT7ls3UECLcIWPa9QzZIyeJvKb
oj+NAIUGlAPZImxbbSfpSjyj/bAcYARKJX9MIxSPUDv9KV+PZhP/DA+WX8dNHi4s1EGegEvPk9Uj
x7x2Xb3ywjKeyU0lzW/JdoybauuJHUdbfw85vV9tUhYl4iV6bR9XDjz71RkyJQDtJHG1YAh/WLD9
nUgcdfImlkMZJo/bJ/4vVOSdFqmw0bcHOr7YEaN2kR8XJcJ7t3RE0Ffab+DKmFblDNq7Z2z0i8eK
BerXbRqOrKzHyXqefa8p4z5AAgqKNMwNjO+x7AWLC5zXhk6stveAdHi5J6jyrgLvIvXWWMGaQaLL
u2A6oqRMjrbI6mroUBHW9Df7lrwrmBdocp8BHajKKYUtxGNdRLbRAvpVvGXKl2TV9y2XaqDHBSLb
e5vLu/5y7kw50je8BvzWvoqkv7thGlUqEdtM2gZA6L8Du5Q6EB6yOWOi0JG+fFUnjREZTzunKP/R
76tn76470Cry2pfBJyEoswXbgwN3fjTZXfCf8579NB1In0y7SlVQlP7SMBBQH/J/sC6ENtiMVefq
QQFL6BS4ljTTqVReQOKetK9Q+GiVs73uy5N5wfQ2ifEvJOnnzaXU9MJclp8YGRLElBqC96LE7tE+
QXMMmG87ucOybt7L5QUvEwhXfyJt7NK+eE+oW3dvpfix/FuzXHP2LPuO7ijZd4Oz2qugrdQPc403
22R8CYaEJP5zz1CefgzV2gIno7dGqnzc4AGNJtJ9ym5Gm4v2an7hnvXIveDDs+2s+rDcSpTroJHq
XiICGYhGK3CtkheNEZa91W+bvIR+8lssc2Kx+HHp5N35WWJFF4UrUXHqehd7SS/qH/nb/xdEEakP
lysXFj6D9yhXsBQ2mhfEipy8vWrY/FtYYRZUCJJhH2JxobhD6yl7HuEocoiJrGvLhmUrUeamkmu8
kcD+bfpOy467W+ObcNNwNeEcx8UrSPmQTOdytQd+v40pCQ3UPrBpseip/ilX5G9U/hlw04zbM4Mt
ODpQ90F4VFgvFjraMnaYB4NYiztD7UJBGfzaNsz8p9+Q/Ux0GEzGuNSOCSZ5msazgHxwyfu/vgcn
+at76AH88XqhYzIMU1w8XlcM6W2q35LB0cmO9ob7DnvCkS3giOjltkAMHRy1ejpaH23pR0XDihMc
cpzy5/lN/pmkrTIAN8yEpurKvPHO7/r/ALJm5HBTIjDbsVNSf9Kklfi5gLpv9gZLQjDGbjjYWK4j
8/jdr9sRpglnCQYeWqbgtnLLOz5KkOe+dUb45H7GJdcNYMjyluHQyePI8n8L5UEIbB+QROZnhwYB
hWxus39zt+Vi/KGW4oGiI5gvUI6Cml7sFWb26YWZKHGmvpLbsogB77s3m8aZcfMa+cA8ZKwdfOXC
JwF9XbgyUJHvYSvbvaXAtPjRCH+EOHK+3ktUIcgFb47FMs4qxK9BBar5zO24+21I1iiQ1gbDGtGb
ZoRB6rVyI5d3llrhDpD62sV5h83PLc7j39GDsXHFQ86Oi67AH6iUyIrkQwEiUrIgtSQpCI9plVIH
tOfcEb64BHwrLEAgC/3/kBhwaM3TOCBwKKJYvJQT/HBpyzMiFSOjY6y6AniYBwOu1JZ5eW0xcGx4
V9qbHW8+vEzZp/3NPnuEYM+erQUR27BZu21sm4WcNtzOrU3IRSqjqVq8iKXWvFopK2r6SvNxjuUS
YkjqMv+M8km5CFG4BtyDE9E4U7xmsBQb43MNUhJa1wdJjgNYLiSqiAUksFtLZ3qNaT1zIoRpFcem
NwDLu6Kp3G0AvCPA3nY2qRYb24Ytp/meAX7SpSJ6JS/XWXsaN0bcME4Js+34clKVZ7taNlhsXrct
7BvpEuJRgGibajmS25tSzdfpveryHXq3pO3eFpjTSZa3Pn///I2T85/F6A0AF7Z69o+EBKpC5crR
q2kwgni9Vip0AhSNlT2iTPEuoVqXNWJc/xfcG437E2xshotfD7UzfG9kf/snt1fCitVOp+whxjhQ
BZUstKACQSVlXd1wj+voYqrgfGCGa7wXCEgt44loOyZqvimvgmBrpCC+dSpKTGw0W1GnbK6I8Dys
viWzBp13rbZ4WjJUzEPIQwpT1bGnMcj4tfsdLSdbF7Buk0LpLNVhrijQO5ucaFbrhH2sMtjCMij0
F7+44Pq1eXkkRV5RbEaM5xTvo4WLZa2B5Z4C6qiCVhwGGG1G82Qkq2cXEI3QPsG6mRSqzkTN0Thx
XeTTxeAIZ/u9tm0n0kZ8XGrjuNhpxAoKgBZc0x1IvXZb2Agfiy9ZeQjhkqQfdwrVhBpANPav2gOb
XvG+LAh/f6EpEPgNMd5p1/G21Q2xgTehIPwHSO9c+Kj8FmOv0iSDhzR3Z6snrnhPrSqJ+95p7F4H
ml391pL2ozZf5NKvffNHlu6VVhlG7B4Ej8m3SdtFuQm19NfzVyTNNnnaPnNlsO64+OT5axig1QfG
AyIHeM+KPa8b4lndUwHoGj+5T5E2OX0xZ5iLKK9G4PkTuLQ5G6Q9q+pcu3Sak6sB915z9AC6dvU+
egNnkko5zlfuhpMRYlHTADQ83+2WxPwr9434htCZj3NST/e/hXweJl+POPjdL8ClRtSUtWFaSKAA
1m9TKKfwv1vMgF7d0sBUcFtTCLmbwUfz1gfOmwVAzJQjSKsK9gpIv2x9eHBIddzlxWi9Rpvds/xr
t3LuV9I36tQ5qdlI0waYbSzhYXQnTmRNg1aqVqLv4toc8lwQe55XCMIpb/5g1uQybtrEjybK+cli
cAMTJL6vLDTuiLXOLrt/G3rPWoaBMqb+LPknNjYb89D+RQK7/cLEd8M+jG1r17fMHodRSshTrMVG
R5Qlq13Dz1Nv15nu2GRtAWP/eJV6ImOoiV9QQXd0jTLV2UQBUzvI6MQRA+12AQlOvj7X2ysdmRfP
DlkSeaq7EO4bjUKe7ICDlR8VA20+tdk7Fs0q0Kqp0v8VyT/1E5bGm1HA3j5uPi9vK3enZCcpfa9P
ZYTsuXoWsfyF0+DVk4upOKnbUww8b48qm2pbD8YZ927M3mHzrOYJCWDk3uUrCr6MryPTwgMRlbXT
dx0/xBYmSJuRxdFdvjcNb6T3cIzl8QPZUajMldcY1tlo81eoB4lIQVIvnyEiC4DVbdK34EY8DhIW
W1KUV1FBPa9hYoRsPjdqiBgmi79SCU2qUA5jCQbVJ2xiyVplfMLDNufE8uVXEoJzAs3Csxl718e+
vb5509fdqvnRDK6KdjujWf6Lg6MCzbrRe5ZrlLI4BcNDRsJ+AW/wYWHHc7SEWV7lQwx9xKPPohUY
Qy+JTr+0F8DlRWCJ0omKLSeSpA+njLZ6aaOmJ2eIdkftm2TjQgwYeT/utylpmvVvVTzwFMsSh8cr
zdIRPb5TdrCNz2JNCcpns9X+CBTRf0dyFn19XTSrIg/+URYfE678NlnwlXeSm/jcecSUNyFMKmP6
/cE/jhZ2gjtDshuLmu+PUS1n3p8hGzAtkXENKfoOslTzXIbKhFDcOTYoU3DBJmyYkAgjZ/B15Gi4
f6z61ixPL1dtpXAA6QPIzDT71TVqtw9rx1uSwBVOw1a9g4zwYXzO3Ah0+SaUkU4i/7wg+XvAgbpm
Tsyfe9R9Ox5VUTumiFM5QwakoomyGE4SBXI6bWXYjrsLQyzHpSq19B04ftJfl+ZzE1ONZkpRlDOv
pjF++U5eknKeHdPrrcqDvdZ0eSFA8HaPI7HOtrNw+qyqKTw9nHF4eJKm5WIm6mZr9YKGV1eC5ugM
JUhBJNYv67oV1AZKWzAkDiDnM2doH5eJUbvbQMASll3gv/rfwgfqFyGAKOZoTKX76ApQYkUvTMr1
xuUqTwXJhLQnkQUEqc3PuWetladmlI1LwZXMq9CKGDfTnb2lPT64O6W8Qdf2+nanN32VZHvqDEzP
RBuSaDZnUxD//Orle49NOd+qqd8uP9uJNOhHUZ1NcOufgvKZb/41OH04+9Jzj+0rJv8ihy6AUk6F
8JYyLbJSGo02z62PeA1GNX43/Yo9Wbb/yNpCwMC7GUhSjFFZ6+4ynuKX0xWGBJzmULuuKFC2hM7r
/hDTspMjkAWiBxTrQW8s4pqgWiGD4CgokFsTqmGV2U7s+7qo/geAqyHImbzml39eXVBCjRbM45KW
i7i6hywe/eRHSk3TWNCuWLie/Hm+RrOw4YBgRpiu2MkcCgt5QiKCYKtdfKI3NAYAJquojdb3MtmF
0JeFqTpgGAcwXvYSixQiYUnCnHTyUpv8PS0eJ/n1Pqvx+XSBBiBIBBNPNMOMW0+bepreb6l/zuXt
uPdKVAQ04j23/UK71nRZN89THE6AbSWoRduc2IaH5ocJhBnfTF7X2e+7wsUPze6215gaXrQUrAVR
uzZSKt7UZZ5sPvdXE2Zy9LjaoIPjMOe1XgL7dEl9Z1kOZfQmoaO+zJ4sRSCLuLcp/MOjddi132mZ
vfYD1T4HJXf2EnRtpAZkRYHIAinZPiQSSpd8IQMOVxStTV/2LIVp5Ixw/aEN8mJUJlA3/0I3Bv0t
z7xPAHM9KnC8XKMxfR8BTr0n1o+ReGXNmIYMkTIV2QgAhMbPtLMi90ZkOaZxZEDMB//DtETThK65
p5GjrQdTLdkHGpbIVem04+8aul9BnARMhziPPwBWDfMtUhlrxqoxPZYEIqMvSfWKmfLMLRyiLZQ+
MXUjG4OeCKnVR/CeGSoRgO3i4L0aLUIX+NNdldn4Cbjd9SYxOedhdRjoGuqo8fHO3y+wvaIHtzTz
QN06iOnZGR92CQwVFQxNVpqh67GL3cBKncKmMyzsBrq9cvy8mfOKdYfkJkK2R/6CItV2taf9aibd
+zX6VJ5nAfjzQ/Eygj0jVHaDUwd/rzxrIANoziNVwg40KTs0h/kohWn8V29fwH1UlmR3mwXKC5Le
brsJnYcZDxS43VVSDzCE1s0gFaXg+qL/EWwnROLTYMdEKZGnWuPKTb6/bag+5veDRNqJDMscWPuU
Spg0hOLfBaERB/FX3nKtRjXShVjMED33wPX7rupyXdlDxJTOatAS6jxUA1w16QBo4jMR3BYXzcle
Prjjk81DO9QVXGqlzNPkiVPGQFyPedubLksgcT/1vbJIUDe2INnUanuRorI0gAR03yRy8UxnGnBq
WTZsaHI/OZQrMiLNtyuIMOR23HJ9buHaJbXhYRwqBLuB1eIHtelPQuX6z/rssTALngsvMwjHyASu
+dx9tvwV4oY/XrtYIrIWRO7ZMnmFLAid7AjOOUWm++F2Kq0f/50dQa/2cw3Te2BiO+rQpWuLVBfa
fao7qVHEzpEpjazZYv3mBzQgvfiR+BnNmAOP93tu201F9YBrzpSmm0tXNrF++nzTC0cKCLXKZNpl
op6Cg8hyjhwzWDS6fKUQYsb6n3Z+6g9YS/BwaafZplQvtE3XfVfigfAMxqr096FjSE+PzI0EV5UC
AtfFUtfIkZmwq70/zTokpEK500lM8NUL4Q1EjYkTJl3FNCD45VXlxlz/0dCJ5w5TndzSskt9AB6d
Z9pZtPyqS3svTnt6tEyUfEbckoFJ/6Kj5iL2+e2Q7//mpfrE9d1pMUasNLVbT2bqvWKq5JOBqAiH
qa7Jw9hxNSZLU6aT4jJ/Bh7AkwhBnnyyj0jzwJGS0hfePAJmMjOTPwQhzBz4nJgEbMglnilwjphC
FDBdDw5LLfdCPA+I2rS2TCWvxzjG6Y+s+dTvjsYlYgRO1KSAg9LBupu3QkTmoTFKpeeoKSuWZZlF
WTYTT3wEHh5jI3qnyLPoAetiu0Crua9AzbhSYyqCBhu7KDChhHJ4CIJycEfPWl+wjBYo95LY/VxG
kS8qnfitmKWUPM2463Ymtu7srVIatj3o/YwfDExEe9YSRPpd+/LkCj2J0Hj9hyzteFNPqEXOebeB
OlldcPPu2Q3dlFbjuR+y1y+EPcHj1/INYP0AFSSVpIfvio5zkCdHSK7owdANWaVwAXTlH3OrU33V
9jNPk+nHU3SD422+7TX7D+Sx5QPnB3QNBFAQbR7O+Ktuax3cw05R6ZJvC5YVJ13M6263tFisMsWm
I4a4iog0UYf4/DVP84/hJ1qmDSzk611A6Uk+C5XL6CM7++ib/4XpUJjJg+EDUCVlDlWqdfh04gBg
uh4/jMbSCT7ffIwCCmjwQ4eJ7MDlRAfehk6v4D4hNXyPdKscvOF6pVF8KiO4kO80YSF8TcUb+SqT
rc6vspqcUtgA+GoRJOkqgGBkfjMpO9onprRwJmQDvvA4MFFb6g32nfIQdBS8fuNEb05oJtX+7xJz
utdv7JMGTDTSYv2KlZ7Kh6nPtirN9fE5Kuugq0wYbVOpoxOb/TzAMrX3LJlE5iBtGatsZdhvODAC
MP7ppOxzaEOA9aHrA1Eatfkg4cKITMRnBpLb4pnKulQvrY/qBvBPa4EO+uxQ+//uszIYdlQ8xatg
Kv+biEivDHU6FYROZsKP90gndmKVDowsYItf/PhtLS7+wE1VpXYN6QkggXiKrwPH2byqllyxqgHb
zp7TN2FaAo1uuAyFyqdWRnCEicYeqKO8VC6AIKoyyzBh52/7MgXfGXtoA+W1Rzne0S05wzIRABYD
g+1RtuKQ58tHTsXDCjd+clmjD30Mx2u2jRApP73OoC6UG8s5h8FC+Qs9HZ0n5dcG+2SEc4Xagi/N
TaBqN+2j0yTcYF19tipYBNQrJzAFraPx1ikZrDkKz4/z9rb+eQW//Iz2qQXb4NvUJlQh87xKU9wp
rZELjHQGZsIzEGR+LnZjenb6j4+dI21qdd5olTrS43nKYPda1HzQalTpBcKKycCkGUUQ2jiFWbJY
7immQZynrgLF3orfFjslO8/hYBEAoN2/ZVcx8ptyE/BaDUOjW1RC7yFFlT3GsSjjS1SAPe+LwLeH
QX1cWiXJgZM8YwbUE2hw4mJ2pxard+8bTAWts2QyvZEzJ7PLuGAi3WdFJFirc+LfDrAvXaVevbvs
Pstj8BZuVBovA1R+sRLqtkLwAPKOAxpkhO8Zj+r4hssLE8FCVpPlr9DicOsdGsiZTWJPvMeurTUt
SOqI1BNqEnXG5v1Z5Cu8jxXyGFmK2m2REFtcT/Mdy3gMkflue33eiL9UTJOXDapb93e7t11H8Tcw
cMyJ9B7+8wjpfZQ6cwzqnVWefUF1lTcP/nD6dzYR4QzaM1lqGDltgS7ixZScDMCR7ehEkXjZxVdA
scYNkMw8e0NVNHH/L5vwwE4PkxdTHrLRH6AFu3wnbn1JM/4diLvBsU76im0/MAwSucZfh6yjaYOX
vlDWp2XXElX5MuFN4EjLnT5yajfVPbvEMVn9v69W9vMgYTw8OmDsiRMDI+AcPXKCiVMiCCTVz79l
436GXXy+iN8VmykDH/1AziemtlymJlYkFpmqTX1DZrbFVHyC0ugIt3OmaKsEqiUsiDtKvTYDar+j
Bg6L2b6aSgX4E2PIyzaallaSGZDzEi+mVJz+ZbuLb837u8Me2P+tltZw//uKlGhXu7BKyC1WBymG
xwYzKzyY480grkNm6pNZLsLqnExXXCG/d4WDfXC6crtaToEVumiwQGWTD0+9EBNLX9uM33Z3Jaxa
+27gYgmKgCoS0XOBTV8L0ybNgt2Xz74k2z++UiNUxuaXM3iSVcyJQPABhXgxTIXX/YVGCO9udvZx
mul4z2tr5Oqgyonm5rHZc7LtCEYxgJHCIXrav/aiX4EFTQtD6IEP1rzfH7tkw9z0fgYWLihDuIZj
zdBb3W14VNpYmnflSc2BKBdcya7WJL4xHB+4+V0CIERBrHUV23UoG95+6RT5ISAHGa8DpqHugWXT
zRH9dNksbeRPDEFOU7LxwhAENG+zoqI8K1EYH430/t1tTDDzPoWI10LvIaSUGMyRbaNyB4titcTM
OAB/iol2ssnGMBd+XmrS1YA2GPwuI5Vrc4uUDXI7dTcSpwcVDolnXAus+lBZlJEdw0C3G9tMe7SD
RRg70m46VpOCnKrRtefcu//8ovGMBwsCwB+MPXD/55B2ERBFqIPy75RdSP6fVw6SghXXeIpgQC91
aGG6m1xfdn4+xnDABrjAsJR0vBUW7868fdAOPbs/e3jSKoMnQNXlfbvG8SJlziPDsK0nLzYFriqr
uD7R6v4qGvPAcSudkfRtbwA/Y1k4OI6ggM+KLgWznKdgIINXQ0g8b2I/aHElZ3+VWVBYq5GjCjjo
LxFIUjR/K2JNY8I7InNCv2YuH+w/r/iNEVJ0lzuLxYHOjW2N3KL/2Yb7rI8RS+JJSLW6VFeGkaUO
YXOD2RfP1DSP0tC8LJZXz8CR7sR3n2nHrfNSw7rb+vz63yZ0Cx4x1VJ4mcp/HzyfWiqAObCQPHZT
fJo4jniOmWodyORZKgmZb/6YN8dgU04kdOYMQMCvXLSOBcnDFa82Ry4t+mzmBsSwWC8p1FUzyVgi
q6BNYch5ZV3EgxoQhY5FsPM6M0DQi/VEiIzVnQY6QWMyao33n2IOICrHBYbQ8zMU5CSjM6vq/un5
kO7D93LPnt1W7lIQ3mwUOqKQwOxMuO77B0nwCkfKHgQnA8jmwk50mx8f9Tfam+r8P+yldCeD0Fn/
tbqHiS17o+hYug+nfslqNkSthMbJILV+LV7kBhkbCyIvwV+LUAWGUOTwIxtGKQ/aI0QUqVRhs8VW
949ypb2c75n4+xSue68KrGH4r0RkydJArHsz1Vc2Ako9hy+QrKb+WLoD+Sq6HagfIl5iROLK62pE
99EKw6lQdPAjMRbJ219Qjdz0DDZwuEo58U1XR1yCfJpabwStwrAGppc061ne8Bls8O51w+uA2vdz
RlqdiNw6im/3MatmrO5GIdpk6m52F12y25blIwa2k1qauNf3B/OhbGJ9WZFnBAtALkZH0tm8oa8X
ItUM+fOMDAnfRug+xanPtiqe0imgF30Hzx5/oMCF2MprJWNQERqwRPzXA0xzl7auiKbkuLIB2/uy
hbGcuHXMaOfDevHg7qFAIqVvdESCf8gn7fVA8E3JykWGaRdVMBFRy+E1EwGIeKaILKF48ciDx4ZF
QtuOYPx7ldZKcpyZmG6SM6xVSx0tlqpCDI1b9q2/C9tVs42ntu9w0Vps4icmXnpETOnxXnBRUzHg
CI0zX/MkhqAF0CHObh0zi+8NwdFtlJA9RFzO3NWZiXgCFrZQQTw0uqEG3LjiLZqO7qtDIpqcY1zF
/KC3O2fP62fS88hIwhxzKZE+k6Ktz4JVrlIjB8oEoWbRkj/MBsCWpO2CXgm5HN3Se6Eb16RYLCNp
wm+DASPS978pIKF55vZ3JnbIOZ0QH7FUVyi5wKZzS/xVzy/tRq9XrXFAPVcma02GIANN69XK/I8F
OfKLpZ5QmfIUbLJ6/XaZgcdHNhYjxC6cFNic/QwoOKNCOvP00hkvmsqQTNe76woFiMZaDwsfLsJq
dVU8kc9M+a+vYVKMk79lwuBwEnsH65l9GIJDV8Io91E3mVBiFP2AgSxOjnH4rAdmNUzlwJXWckXn
2Y6zYY2I7s+2+Dp/QCLCppPYZxrT6LCbCi79lpivsZ8GfNW0qFmmC3ociWlVbtL17PE3ysmAE9xg
arokb4vf/EvNasZMmFoOUM9dtIS+yV5szNDRhyLFFqX+eQd6/dAp3m85Fm2u/7IUQ24OdwT7ZCbW
NxvbGZFhGo0Hu4He5X/OY2D2LjlO4Ga0SkenlY3vTPKmMEhDCq2ZHpV8gFzBHUc8uiXnlgXh27gW
cWi/roCeCCUELLbeyCFeHcBL2sWhZjc+2yYPsWS9T5EMQO2I8vYnFILlZW2KaDDyuyAiCD0TrbUn
07sYJXrF9qxpkkdXYSdO+0p3mgtTKik0nojI80W6UJjt8aTBk3eNFMLoYSQXuWOopqRjqnV0kgK7
lXB7jB83aFRr7tW+pNLk61SisgaRTS3hOLKwXdQwo1SYs5HbD8MXKT43ZlUjG4DV81CseeWClsQA
+6nvMP/OCidnvqnQlHYchJjbLwqDGFKR7wBS1I7f4pqVne3PERnDUZUnnAZBXB5hiSBemux0hhN9
WjmbgtnGiLN3ZviMCvXU28HexCWUv3cLPOksLQsEIZ65irhfSFul3pmSuhmVOwYHKZJELqtCpQnP
PnmCPsT4XL+7yyNfnKiU8K2q+cy8YDzoZanD4BhTSaHaNWHNWS/8ZPepweBIREoFwNoEyhnN0B5K
n5jHnghifv9fURRzujOxJYwVAh5xUX9+9FVsRVk6lFToacqp1e5uIH6HLPPtqK21aLuPajReWeU0
p1Y1ZLtuWwI+wJ5H8VfgnlIxqVtEgoplwO/nJ/zjQDfnnXfpvKiUXRT7zhj0I80Z8vheA2kFSHaf
OAkNAOmV4BuPq4evf2+OYc9i7NbyRCvVXzgLGpN+gta0f0j12vKNVsB6VHul2ThJ3Izx6gY8yWea
+PaiU/TSZ0F73ZdJRUDUV7mqt0BvHBMhpx8+2DZupmEKv92QXJo7JSEVxhlNgFwHl/hbVPkHE8vV
2wKpb5eT0Wvrj0iG84m5vdYIGlay7vAjcAmsUcML/LmV4yWDg2Q/mccWVbQWqZiefsbFsAve+ctT
mYDqo3hiPgrVJNYSuf+mKhsS/yYers11Q5PljQBEkl0nknbO+9NkM0ApoLYuXtJ2hs8tkLjtNQ0s
BmNbtMt9i+pjCVYBSYS3JZT46JXUFzRfNCWv4n/fwE5lKeRbX4tJ52oyC5pfKYc7wGrTSP2p6upF
iBPuhKKtHeheFb5SQqWtaY1Ru8rkbbFVNa9/Y7KdN/xwZR8FSLL2Q14LDx7Fe823a9gHsnEpd4Tj
LAz9WajlpTbLT1MbszWhDKM1dO+1A0QGu3uRIfQWqzhWy9yf02Hu4Bqek+aWdS/ydJW92fWbhrCH
G7Xlhn6Gm1aZF2gSvuQo5B+Zr+9s0CS4ZFpK0eJ6QYNCiOebKwysBlrDKFVD5sjdYBiaysS0OLxR
vj4exRB74yZWPr0kx8ixGzJgilsVipljwqQWW6BuM/f1poe+RGgdSpuAPiqwYzP7VFZZ9x9MAi4b
P092jto8g7e1ki8ghfQY7JfFZuu0eSPG3OIuNyk7E+RkVM8D/nxGpeU/+RGbhIgq1XVfHbmiL2w2
+TrsjUX6It9FkeHg3ehMk3bNbhh2va3gaXePjH15IumsoFH/rLirT/w8d5ECVZUtX/6grNFb+9wN
Gtd4WKhsCsDuoxfX2Yn5fG3yr3qMcObeJPrT7fn0EG21seqK7xu3s1KO4ox+P1E1s0pBeRDkHJ1X
J1NFHTpwS+WZfy1+zVfAbsK2+UO7Imui6KMm/yBzc5VrQP/cbKAk295f7P9ekWeEp7PCcjK8Lbpu
O4tTU9/nTA20j3f2E00uNVk89nn0ZanU1y8ChzFKyLwFTTBe5MTDivdo9bfeU2lD1ppU9Dbiwl4K
TgkDVDpA2ogbRIYGZeN2QZRPtYarslbHKe4I/XlmeMxTLY6xSchKQ0f4RlrlfsNU62ae5XdBMJu/
9c+jBJIdVZiaVzdDhTq8aAJ7Apyh5RB+mcuFG9PnUyNwWMM4uhlfwAWY7p9Skhkc/6NMwhJSRk3F
tMoIADb8BFIy6zXcM3WZ8gxHEHjLMTzUZbzc/FgLpp0+9xG2xkwTWa93K0BGvh9au6IfmVqNheDw
ubo7pGb2M+C66r9vh2ojR5Z1zslsbhZSImyy22uznFtpJctoZcLu6NRMgFwdCfNJNuQyqOMVawIA
6RyzfOndgSBZWYu/ezcK0F9xjewhEsUlNYSK8puTybUjQzWDEIDYlEzo6vgOzCnXSEYABI8Y67Qg
QVbStqLFZVQcTF8OAVxJffEhd/ZRUv/HYTJ/qtQNhZFF0hc2GkM9ZyakodCudBdyZokXxO9ZjwTy
o7VWNvAlB9dN33Y4xJwN6YJMj9sr3WwyMqwJR//0ISC55zAVY+MXq22qfbLczI6hbklJFJWzsLPK
EJeNQhuCHxd/bvUZuJ8nCejHrAEOOUDrz+UUN7rv3o7iaz34Is8Skurik/S83MAaGpfbuAeG4rZW
THieq+1mXo/sXegXx66daK9Pvv+tLfDQPKIs4tEooip/gO8L3OdSaO489ICcyO5E2+Ve7NhtfeQN
A9tf9L32fC/L6UL6VJQcbw7ezD2RLKt9azZ3o49mIZN9O9fUExmSredFd9iGx4Sze/CaPsCVAOcT
hWTRWHWkUcpVFpL1thgRI90A9guSA0TDrefG3Ua/r/YkShsvLCoa8BbDyTOGBUOSSNTDDQF1bt/m
S7k/Do31FXbJQCu5ZMsmVUvo4qiiy/Zl6W5MbVGuzd5lwQFJj8aLnrCnlF5oh07ysChXTi4Y6Ppn
138gg0VT3C29Pwab70u4jWNVLcbNT+hWigi3bHahAna3Ru5f58fUwabA5GnIXRcAsjmJSttHSC13
rMtnSsG5E1D0c8oVIj3YduKF2c3ORufYFOarvXHK5NV5PkixESSOguTWEEfAEolYGr1UZBEltfsr
kY+51j2qXZ7P6lDJxgoZUquossHK7hr/gmsl4XL8m6kGezQ6Wtq2pqj4SVDLveZ6SjKJUzVvSQzX
oE6fW0HkiIESd7mjh5PL5vdJqpuD87TXlM9z5b3U3KvTpyxvaDdX92ccBIsPV6GG6hAJdAloEuwl
7kd+9ypdcbx+ftJbu1KhngVpQLSXr7b3VAqpn2nbiFm2crzfrHbKYUkI5dz18fD7n+2Bh6xNB0oy
vEl3uQDxaEm61CVuAJZ225Na6cCifHUnhSjyt6fDAGTye5bv/npRCuzF1FUcLhCBXflC1sC4g+r0
qtzXIqsUl74soJyFovscI3hA7FxG3WMymaXOms7gZFg3E4yLzRs5j1pGxzSRJ3smMfSBJ9ylRMCd
yfY8bB3xPNOxAAj2m2BtlrMnYgUZEYDYkTz1xy70mlndT6BCHRibvRsJ1FdVZ1fZPjDboDUe5bK+
aIdw48KZE5TtDVNTGlgeC/MuCeYGFdZgQsZEsqEjZELPyxXTRzn9yGMDXbYILRXiCu9oY/IEHbj8
BoCopIcwrG3z5/W0AwcUPg6ORxRGnXHucDQvDfUdSM56oCnuZDaa3d3UkL+dTPNE3gvaFX//EnBl
9j9tQFoQD7MM2ral3RUv83TzJ5RLxRoCmE2LIA4JXXC1uVWlShSIBPAqNvO3YBtOUPPa5Ujf/Lxy
bhJkd8ywybdfKEIXtxITFDUZaXgtR7AF5ZaCAtLN/CexBsf5yRFcJ0AkMOfC8/DgxlawLSXUbQvY
yTH2YIUxPI8f7lpXrc22w48Ti1J/OVhKxtAj2N3Ukp7MBbnM9DvhGEcFSIzHJxH+PGX8rh0bP+cg
sr8ojWrFoG0ItFwGQEqd+xiK1Al0vFXPUtdPHOxfemnZTdMuGhHDtX/n71m5Cub2qSoiQA1p20bi
sxmld8HaJJ6VFMhMhfEZfAPUhse6uacjJ/ellIuQ9rMmGl9ZMK49TuMTlOKzU+kQl/mmnMZpHOEL
7lcLM63yzcMOHLGbVZkBqC5RiV88609CEho9X7RdByb4pdvLHZnh16IiRjDjGJF4cL1QfmcFXqyg
joAI8c0oWfM53szWXOf8uPssDGc9ZankTuGO1lxIaOPmeizlehhKk/+yD1kZHKG9X4um/y/uUjEM
7uX55ESAe5L/n2tKvlI0MUQcEqpbxPqw7HJZLUVobbCbcpF6SZAQichzJZXw7B/EzRX9UgJeuD+9
fuf2Zgsjp5zMrZB24avW6XQ29sK+RVLA0tggUHN1woAdDH2MFIr05yXVHY+eyZnrpvoY69T25GJL
zl/4vfR/4gm/LfnS3SDrk+pBaBfZEoh87xjTuhv0nhumZi2bL9/xnDDYk8gbsH7TKLRXjYtB1w2M
VgNtXRc4vJCVQz2L6pGUb3xiOt9h7bNK8ua9EUFvin+Z7UYgduSap/CMY0sA5XRrDlaL+Y4ZsLpY
XV9wyQMq3ztV0+wBNW9fk8RC/XX4ja6PWjLvoR4DlLerAkQpObZLaxwQvUMNvoIB81l2DMpF54/V
WysXOLIp6vDJPTaWHwVO/0zh23EsNQNeAqyXI6eTZkCqfYhDTx2L4HwJwbxRDUGNfwRKMHVLQfVF
f3IWKxolDZCk2PNHqspz54Awrdu2FRkZY9ldXkNp9kMtzVLJqt474UOJGjYcsyz9nq5pfe6GRJbW
R1abasNflwEXdqunPIJ4UkoLTahwVu9wNnSeWbwmcKCsh9HnaxnaT5fO8JbqeumipaFjS1mr6Npl
jwYIU1SCsKRNlLS1n69mBY5VnkPx3+uyzK5CoS8v+F7ZhyourpotviDYmwUBy88/C9c/9dPW1QMf
5GTIPCMAphyrVtLP7j4RwdEYAOJVd0DnHBSi08whtyBhQXSKYmPLm6iEwSdpbHZhJmNfFjr0UnNO
t83wCpLCMPUGXzAWCG08vWqRnhTBuSF/rZHSqp+OcXf/PV0bYkY9vSDs6apBGKu5oHt5aNRKQFZR
p8PybH6Lk67hqn/Piwhy92mkNi3S8HejH7nzle3ML6ldDSnSkNVI3W7UmMlvJDjrcIaKPrIC9s8c
a98mISbtKRrjLA2DFxJeZH7gUPyg+wHIVtzyENUJoXGTxKsHv4utZbbFGvUE9KDLzYtNeC9NifCQ
OvHTBgVZ/vnmP558DMEezHZZzm5h/XHvlWWFilgmXkZNpBoPwSRWxpTw0Vi0UTkMgUOSheq8Z4m0
Yww9JH2lhhz9fGlifPegJwPdOmQyCw58gDTG2J38+Fdfi53k3pmideUxkK7b2bZSgGEIqcr0GOtu
xFuY9Bv1mRMFZZL+JaugsoiBo3HppcGNgNQT7HdTNT0JFOV3ijbNxjTVZltbXwSkkCL3EIlCHimY
qt3lEgVOu5m54W4zGcCwwVBtprC8W6HzOo+7+GDmXPSFU97PgQrZ8c3jf8ZMtIF7uJEMI0G6sH2U
e8Iwj0UnxQBa06Eqwybo971gBdNMFkYwOOJYYtdlinLxUIU/zqtGbE9oVHl3N68K4r6uA1H2u17I
Us1bj0JJ8aRUs8CHCt6CFAddynm6pQjcnSp0NQ05rKU8gAjcbA18kvd/2mU8gLE/KlwRvX6csMmM
16pkDxdqp1XIoe+3agdIZAFF+Wo6jV2A8jBMWSv8pWyMPS48veAXic1RjJd+cVePlPzuFVL5Fo0W
b2jj7V0SHWiOihP6oSji/by31v1ObHQlxrPaipEjuuyoB7rw2JFQ5BdTVXFUCA5FLbRCKp1TDr2A
fgbOW/VvCRbNsJ2pumRA9YbT6AWOiPBIoFjNglVrJQg/M/+SYcShMesFKI5XgIdtQdHJrCdSBYk6
7Jirb/nD2GR5m2vaL4kRZqob0U06AQwjzOHj0lebv0COgwrM/fGkagUA6oG4OTXFAd62AH000wDE
JA7DCtQjbMAVVFUg6iboYJIUAOv5g3LZ1/AuzauV3MwllVkjD7Kt/H6YA1DcnYrfqA/fL3zOyXn0
9umjyarjmWeCx/HOTCA73TngxvMXOxkUq2wFN0zU3Gq0iGLXKMu6g22e2/gzMaNf7AWqr99pHKAx
FjmMgau9uYy0ttLnM4mNlt7DxFbwffFKhF9ZGFIx7XZQqlBPzLMuKPf8x9c/nJQdNuBUzTg+Xuzk
Ese41YL2PpVNCi2ppw+9fF4iVAXOxGHirkpV13YnP3pq0ETx3CsQq108dGEny5b8SqK25ESYPSdJ
Cm5yt66mvlM5HU2D+GI1TmSGIroRlQdiYWYWYzBTmUlAnFocL6EyNjP4PAZbOY1NksyhxThAvHGq
zepg1qi/VSDNv7WiCSbbvQn8EyK19++ECAM1c9DT0/ZtX4WVocQTt2JgRPe4qriG+NGKaVqnav+P
Fwsh/K9goQwwaHXhUdpp/J16lrpqNf/8dRPtkRkjONWz1WB/YCC0GXLI4+mmMBmttNC3SxwHxigM
2i+Ibk4IitmglF/kDTgvQqro4s0afrUcj9JuQMVJaFFSESDY+yU99NChBtsO9qz8qRHtkQb0Vg/3
TehPyPOoX14AZgGDdhPRizDSvP6XPm94UZt7WjtHdRucErwXaOlX0YPeSvc8PVi6UigaGzGZR410
wKuBHzEuBT15f3aTlTf/1kVIu71RJXzaExXGJneEtLxM0ux97TQVlyBYxSPbneTKPZVUrnNjaAim
FYYe0eP6n2yc+GjzMF5XKXq8DEgLCWaZHLvzs1aTDW1JkSKrItbRwYiH8VPwahVDTZgNh3zE45eD
ca0pXdTpDJjs2qKNsJYYpu5enUcPu7PUIpEKe1fzBQFGzjRAVBYMoDSQBuRLLMy012m/3wPRWyyN
eknIjuZzW7RoZpooyaW7kxDKsvW/PsZm8LVpadzUtzDb4wUQohByenrY1VFlsmlndumzSE8+EkUq
rRVxT5ISw74jrxqDbB5ppFWTtQ3P0Cm7s/FRhdb8GgCVDhVOAQvh9yupDvz5oxBrUoC3JnvkJajj
AvuoF0JYNCWZQJfZFouk5+j/khbh6O4AX32CdhcPji62mKZ/5t0aVrBZgPzgfVDoiq7SqP54m6+a
48aWMMj5NFwQrlRN/xRKFP81KyBbgEEo6UiXPL87dWApbrhKzIe+hle2D1nmeR9IaxErE6rFQwUL
6IzwcbIn3X4FY1npyIj68KOpPCUOGyeEAuEtlKEOTNUGOy/w2aDMMkRB7mcgZYTZsupLDv4uU7ZG
nVQe2cJ/59ywt2S8rDB5P5mcC2iwHJhmBKL7cDCqS3PmCl0S3RfwnItlvRUoe4Vz+t7mD9CTOqJS
aaA7h85xX+wW9Sr7NLUZoMQnDG8iamAzM0AkjvDEimEkBtihgk+MjsFs1GLRDihsvmdofQC4pc5E
B/3cCwXzGTMZY+0gT6ffeIhd/zJE4ECx0Uizqb9QgARokMnsByxeZ3Vudg6UL0fjGhahCh1md4DJ
imgfiBGCmL8rIuuBmdGEJGiAnzQ1QqB8t2z1j0W57mZEbdPEjTTwb3S4aSQE/e2l1z1TWn5dvUde
Q9lXtfBTR0+mv8MqxxDEfE1wx6Umidm3xn8D5c8PXqqKAVJB7jNWjaK6yoYjFM3tNbZeGbB7hfUZ
DjSytgIgOsqtwRJbwb0JwjuxdP9qCBzuY4poc9zI0ahKh12bWfEaHRkXFDjjE8XbUnUJ4e3CsXvh
yYWlg0/Fn4jj5iQGio8pbhkOT9DfEtOpv9y88xbQo69iurjeHKg4yu+kh4Iq1Ba0IUKbvNwMnJB9
brwKeQfKqdFX/AGAd8GhEt+tY0ep+zMg9QRn4KhOIh6TOEehCQQW6Q7sG/PAKejIKYHVyOroiY7G
flOim2aEBNb3dXNCyk+t33LNhm+gPEKpOONyQdV0w07uJeiP/t6Fv+ZnwcvjoJ8D2KuvefHxTntH
fNJShLFwrxbmwG112zrhc1j+DYBq6YHoYnLtK0ovvtcsCazk/LDdZkqVYVMf9IAZfR+rKykbhiWc
PNVVuIOtBsIXlKLwir+oDboZC2AWQDoS+Fix0UUVj143WA/M1UyBXTMyq1hKfw+5Ztlw37jQZMbS
TMZVNI+5x4aJo6XbBWS10F/39w/vgE6QnOkOg9nZITT9AyiKPFxjtVa2SpYktAIDCXwMaq30rK1p
sz6Qcv4TC455xP+OBivtlkmUszQjt/BSdm1I5fUQ03iK8/XTQQfs7LVAGBCpn8uJixx2E/97dGU6
VwLrVcc48a5cqqeiclX8AR9KahW6psXEe9/xlvs+vd84M/rSguxLT5IJT4+GqCX6rXtJiGc9DYIO
cTYWlgMMnAJMFH9UtKSfUgBj9MDajbFkUOkDprVbP8gJ8/UICUkj1+FY+dzvAe78uNUAqN6SDJg8
tyDY75hsboOxKwMPfnTsPNpUiA5GwWOLgDL6B6J/4ZyAIlqR5lzwyF1TbsLun1z2LXWhIxrQq/NX
1i8y7+VsyBakBoThUzQU7DZ6lt8DuS/3AA9cdiFmaZFDMWM+kgPKL1JWpj9t0XzZk1FH+bsbuyn8
8V5tv0B/sY7XBpsu6CCX910W40W+ZH3mbGDfLf/QRmNfH3tKWj3LrjHlrnLprj9wZ2eKapI1l7bn
vmP8hao0N74ieeTikPZy+LuiRsjDtVsQceLTV53gUkEcuEi2PtW9/OlTFe+tfzscSuDjiW1mLv/8
ng9exvE1bA+t5B0/NabBBMQPtZM5Cij0et/WN3D1WBgGU1VS2LYZrm1Y2WgOJOPxxyGbkSeVgmkp
U4Nk8J0N045dfyLh6TFkhvdwLn1fA7BcquM0YsIWhj2PvutEVkTKeslBGKdlEosPrkgnupkI5gJv
uOrk9EDNEjrRnjSD0IZcnf1A1sml9rpfacssgcCgxY74Idb+ElhbBmCfD0QT6cjUbI3Nm9AHS4rM
RXPp3AQUfD7IqQ0j/ZgXLbrvu48sHs9JrOCYy/MyHlQuHYaAkzUr3pn3cch94qxvGG5xakL9Fzwy
qBYWnYUD2hkIOGrJwVpfW5L5jTL78O89eD3x+TEOiVAtJmkAPD1N1XIsvw/Sc6NC5c/P4cCUZUsm
F1yPTj5Um+I00T3uZWzi+y5FSVoGVoD5PagKYFVaWl8VUj5FIP7bqLKv/retYMlpUqLllwjq8KB4
IgDsvqvGq+wi0Fs99TDYrNXU7geqepMeSDRmm97L6s6aVLR9I6ozpDKK6KFVIVvtWK/1oYGK/clk
esDfWIWI/CAOuuZsRIZeiBhWx8pRhS1kNH2TUuYQ3LULvPvUlwY+ldxxux3B9OAasM6yDvyOr8Vu
Mxdk1BC0VEFyfyRg4TsCrlWS1dFwXYt/SgREUbapI5HXfWhRSHvJGq+0EjeFDPphwFVooeIpb0Ue
8aj8ejMDyvSJQyp7Ktxynd2PZjOMqSqzF3VQgeWNLTEYuMUwh0HDPKQqgqNx9bB4eoo3oyCHbRBG
noRpbmGIxQan1WWrHwDTVXVYjuDN1asPl0fPJe9nwR6aJPYk/FQ2Bc/3WhhaaxzK6mUQymGZc1fc
LM1uFpeLMVUDIRDYO3SM3xjubCEfYl6zp96c/cvy7tLrjREXprCtQLU5qQwdGLEmxAUh+YMnF2Qi
MyCcFxe3Jga4Zi+EggWHJVgog+64SKAcb1rmnpzkW5vNYDghTSilwZywjotTNtVopC5mgOn5zwr5
sCF5kSv9jCT9DL14+SNq0pOngRsCIzFLclLFS0Ods8wuiMqTm62aB0i5QbkwnyOSHIemGpkXMBPd
0gIYr+CojzoXXyu3xuZ9InzmUBjnpl0XmLqfRIuHmFKrtDh4ghojYg8d1HLdsl/FoTD/dfNI1QVq
QEngnaoQ0g5sXFONDMk0+IobbWQqDDh/clb5AV+KXgq1Ak4DIqZcB885atVJ/tssIK33V654/Vda
5kK7kV0/bn95QXRsOAQl5FqKBOnj07VoO7d61AOld0HNkk8WMnooUO9LcmK7Z+dyMSdBYC1inryr
XRlB2jIzs7w3plJvXFxNwNQQUKIrvJSynTGi1XJPWb6jwK90tieqwq32vpb+kMu5UURwrH3B5Wh4
XuAtwxaBDQDAzXLvUv35Wka2mjv6bhw/Qc9gWDsFO3JAIo7VPKSqxXJVGKPZjdbp2s4olhAMyVMq
tjwS3rgt5oAJp3sifIZ54BsJCIgwQpu306hPX+bCWI8UPAWjlJwW7f8n6CRLeg6GZoMYVzoUL70o
CeL3gDfoVSWw/r3JiyLIvJ/5rWMY/05xowyJbDpKCg0VfGQz7VzQiuBAB00BnyI7aydrKY1Oqlti
zGuv8nXvqvMQSppuonf5DyzSiji7gKM2YNuk/gUFPTD6UCkYCTlXxUpg13ymV70XkU0fwbmB++0R
xtwwPXVNQdcb5r1qQY1ttXiM7i0YR/6pEvhejYlXppVcVt5Q8939lvngSTlrSgnsnlmX5e5VdfA/
l9JgiesFxkw9IjXtrKxqWtbu6/RFH7zRqa8t2Gqz3gKiTxjVwd+XE2FYVJGYWKA24euXKr0tnFD5
2HxCXrGao/kyf4/stNjQWv/Hcs0H4M9TUp49USaH9jbDgCaokUihrAwq0MOSg/op2kutDfk3ep9Z
XOZnNghediA5RROUv5YuF+q+Bb5gq4qqVJf4BaScd7NCuvtjF3UVtZW5gLD9n/TZTNfSqKJzVp4g
k/sXfwQNVKpIRYgt4hRcMYYTdTKfiasKKxfubFELE002mj3EbBcHiIwlBd2SNDVFjJlWh7Z3fO7z
28CnTLYnODEiDYGnPOOO9RrTIcri+X/r6OWrWB7Mb8zk1cgghS3pJZcNGh8LAFfJExL5jZGj76DL
RYHmjHaKKHFqB+vtdGs9dLjKM1smo34dnCIR8dEwEUpwSdv0DdCciqhZanDK4jFYAzRM1KqM2EAp
azjSjJIRZHb/Z4ahtbtM9WcSVXz6AuE1kOHV6TCpXGiR1Hb9quqK0OqtbXy49H0sxKVluPa8g71B
nF/CvKgl6Ck5TqFnxekY6816PJ8om16vs61d2DNzd2bLTGI0dEQocUj/QO3ZBzQ/sqi7N3dc9SVk
kzmD0gLN2BHfV+wWKrxQ52D6dKJJMNpPKp+GkX1JHx57240+wdgkF6DuqtLeHu0b06Kzwr1YtojI
uErJwiWB0r+gtPuUFfPQCIZVLln0glTRDXv46Wxqxa10r6IAnJcyc5L0PlWYm0gJJhX/Z9JF++XL
D+eA6zGatbbznMbgFz2Firof0zBWHygrp9LilMrsdKv9puyarAxX/0FANFtADiJVzIM2I3MDjDaA
MTA7YeO1gvSdLFuLba1ghjn5+agFhp6UHdHhquOD9ecUeKnQVbAgviHdr3dkL/6vOTvoUzryXfOW
KcIZyRuWx4B2Ev8Vvl3veexJw8PSUNER9txlHotpuom0pYMV7b0eh+LBs7TRV4INGo6xqSRh70qh
ye0km+JnLbKO1H4eEr+FCnSnWOma9/PyYuQRpEGhasexY0SBQbwORZZuwC/LGtZSP0MiEfG/Nm+o
okpab4qZZo6kxrU2JqAlWD9dzmNFwxgltWVSChvK6/EqqylnaCibjoVSqQYhCF89YsuxiB8BRjoy
irE8/4uRXuAEcSX/pEG6gq/kuvhYA8XmxkWShbDnTblMNWtKTQ4tKKfn15NqQyVvr2XQ5vmTcwB0
mUeRRTLi6498x3Sxyx2gQrJuYkazLFM7t7RT8MpLG5y+e9UC9a9Ht8hf5Fm+OsfU236zQCNNWKj2
oZzmfvRSXdf+NyriDBehUvloYsbKFmbuRHBF4RI2Qhc19unE0npdVSNY2oRi7YiwENNdFMQq91E0
cCiysFMp9uIA5Kr+n4Q6kaFP2XFjtFfSZL+6SpIgEwAdmxNoBH9D73aoYQCZpvfhwnnjJbWweFK+
nVfWLJOMNqt8RQB/5pjkG9m+q1pZxrKMdJDUhz6fRPEUDBvLRHBW234h+jLF6gIlnMQVJ3Vn71jn
NyKJWoEZ+e221filZcDIA6aym4yUUexmU/nqAn8baOPT1R1YQof4HUrLOlyXEHY63S8qgsnoO99m
QdoQNRO9bcGTn/RCQptcGu9CUsLsidpHxQdBte2dhVZVdI4K2CovMM9plZKtHVjhJ9Y2l+V5NBVw
Uf+Lxe1lwdfbrCi/X1158TILp+e3Hq4XlqX8ymBusbmSgMgq9iX04XVtD/b7adFhesYmNRhT4dZl
guGLUge2evj3Ps76kF0liKzt80/hD6GAmhOh5stGWsaDyVXwVLUQ3RsWlkl2+BYTI8XmPLSbvkHk
/Bu+hW+x7wWtRBDfwwYl9oD6EMhtElvVTxz7fxNrJxEcwPSKNTZ+nnbWozTM3VezxeobFejEbFIY
c2mTOzc0g3US+GeophisYmSv98nDbpwCNBCucgKMJKRQGQMfEJXAS0GGG2JcJ7WsKLR72VREf4pf
Tszd2nKNfIrJAH+JVST59WFSwB2S2gnV+XRr/E3r9BMO/m0UzyjFDiUZPoZeNfHRVeA2lYa8wDM9
jZWgm6PE/QRiXZiItsIpXfYabZHEfxRLdXgT6fVf466GeLASbMUtjD7Avr44YjNy2QbnDIECMwTV
idYpjewRx+q9i6mDj8tOytf1lZ64cVIpeb7GQ5I5yf0J9+IPmz4DRa9CJQ302KwkJhW62wnxvJ6L
fo/wBNLBoF6erCJqkwSMpGeXaDgY3AT7RmO2G6GxSmbPUWIwAMlKo1ppkIwuWZxiK659LKOXvbt1
NIpH02stLO00/D/2FPya52PiyXV76BF9FmD3sL2NEHf5z8i196Ux1QXXIvxkaeGQ3z19qHWXsBJx
FQxZT7P4mkKKkUaNrsA/7EQZzzZxU/IVcrESmp5XII+HV06QB5rI3gCEs2RKxj4htLEYXmhQdacJ
WaFK02fqvmrriXjuFIYs/ABB6XGRLBgdNXcAkM3hD/DBDsTLYF4kmYK9xrf2wUepEWDqnMnoGzmb
erpSneIxVfgqy79yfvcgO9niASPM/kfr3jc8sopd0uVf/j6hL70J2nIyeLL0tdD6oimvXDr/29z3
f2AHCC4JJL3IncrHkqX+5lPwnfdDXmxJud6arYk7Gsx7jJz44SXbFyXziO1r0lZBMDAVn/JbsWfH
dh03rxp6XyQvInpL7Hk/JlNJImvcrBJB3MfxCjPEz7rkumedQnTkKzuz0R21MKzN51V0KmBvy3rM
8398SVFU64r4kC8HvJLxYYN4pNZF9k/ZFrxE8kQ2km+wV2UrOrGcSsQCTEzailLXz1Kt5piVtsnL
8a9Pe19eExHvPIOyb8L14/nIoEVTPzcwGi1cdKRW6S7P4VKU0DeWBYX0R6+cuhAOgcot5Ue32CgJ
892JQIkIB4BzqU8NRbMyVmekIwV2kJY8ArKutWDEotqqpins64QmwcBNfi/L0sFdjda29g1WPSMq
x5ZUBPStCtE2YkUm1k5EOzgMNWLBiTiV5l4SWgquq7KrXMR5IcO2stPevISxAcbI6NTMY5ahyOap
tp2FE95IvDJEcEnYL5KRHyPhOeWk9s9qw3S99AmvQrRy+mDZa3dNwzMi+upk6Y9bs+HXsiI42uDV
qXqCuJb6kvy82i+aJzsSBgML+blWHXkifHWOXJ2Olax0buxBvU5bNxZAgBWJOBwsK/UTaDQC06LB
7FzXmArwfsrPDg9hCeN9HcnepZoGpD/yf534XYOFkeOQymAEiPWu3Q6nkzkimRQxSNTh+Wnd/krl
EOQ6YA1cERXjKOrVJn93/aJ1XMaVGnxRCVW1OAcvLjidZXMigs0GhuoRu0EtiC5i8tnvOsNct2eW
bhlsITojogdmBpMao8LQSUZ/zxRCkkFpDN6BgcnAqS1B4WRWzhN32Qo/DJ8fvJpIgLU60f6xJbkq
c5kfMXSqS7XqKND+sZF0IhmlB3MmM+DwTNiYVstwCXeGZuImaXL5fdaG6SVSrG9ariEKk5/hD5Di
veP6J8i0A2TBNbxmvmD4Oaehao2SF3DQP7Hnas7gi4HlQW9hzZZaAtqKHyRtwE0VxtyMQJEkjMvZ
H8fbZIXTFxv4fGtXa/3f9YJlS5E1lEc4WLET7eQ8IU3/yRqQ6bn5npjhkxfbPCkr/d8h4EHKcKvV
xOwWqLwvcYPGc/+j4rWFc8MtOFhPHEp1rAJACnlopt75rgxtN9OZC965wRIrofpJ9MquchPsPrY1
TdAiDuZ50lXTkiJol5vLi9L3GdZvGd8r23wcsNDDmic4sr6csECH71NMSIMx3SXzoRw0KTVn2yOA
EGaagsq1NnOq+MptM61qh9vXbFD75aBtLPkLC2dNJ/uqursln8lwE4RtqXFL4Pr7XuhKXDzTDzHt
ihb5Q9jma/AiXLLNLQ5cBK6vi+QVcM5Qei+ARwggpGz8ZHsPMnq/deXYotZxvSQqDHI4c6JKawJv
/IlXG5mohxrbBq2RdYZ12HSMUpqSGVcG/bgVuZf0bTPxjaxjyC49uJnRkyyLmBssu3ev31l6SnkY
pc7PC5nsD/+LUcoz6KOCmTUMJwSFAi/JrMGdNNzJU2WIrXoBWlB/4vXonsbgvMlHcw7I4e0LG3o/
rI8XFMO/35TuEF3Bd9aqSYfMdSTl8QL78CdyoYnFLIWY6sU0djGqPnZjgOLJwj0FYmeGAAKAvas/
YM+1FX09ehq0KJKYXyfY38puJpbx/PGT+szXKkCkxkINehfCSnkDEPLOZVvgqGVxEoWIWnVJDNIF
tUvyNpfHt9Dm85QWm0AvGPcwYqSsM/d6+KjbNvc6R3DTUMczCiIefCWdxIKpbq9qpJ3/hbeN9cpX
1JQN6ZuPqBGoWOnvRofy3r51f5tT0+LtQfAQItvAvatKZz+iMTK9b6P5u6A6bwZXk77ZlqVK3yUc
YyLt1H87/1a/drbgb0hfwwdXufvgOnlF/BDpFqPPO30xRXZb065xLmu8bbPPau9f81Ur6SRBsd37
RDIDyyUQtAPOvX3Olgvi0XT6zRufK/eo9+Y3CfA6Kh5tMEGGP54MYX0cSc6aCRVw7MnUyl91AUYZ
8lPZQher97DEuEMfGQ3WMzEa451gUE90PkP97tPOvfNv8IY/hpbCOciMevsL5cCMpP3Te4Rsu2lk
wGI7FfegEwnPQUZe5laANvBj4l5HPPE9l+DJLFprogCeP5yQDMQk9wRLTSKH55/1TXoD9CSd6Av3
rJumiOXEQkWWTHEpi1bDkRbOTUuwHBYLKYYuc+vGJ9dYmnU/WpNe0JHJiuAoe9+6o6ZaGiukOl4S
f8Ur6wuKk0vXtcwsQLzVF+Uv9fKwbc2TApN5E/5jb0kwYMAUwGOkUbMkaG+Z75JyQP0i96clZws4
sEjxuYD36dS2Waq17DhaXQI6tQRfoX7nsVVFes8anM+c/XrJOR5OAaJu8KXxGTuo8GYoFiOH4U3A
FBU6BBpEysObjMcfuzjpKEMSClw5CDqOid+h8t/1yXtciLAOqhgiyosdHc7M9AHuQXK5MrwJQTt+
1TR14skx4hNCL8qyqu15f3iDbnTxYv6a9sF3rmM28zU9/h+BqeJQwf4vTh16Gh1jpcU7y+3s6w2F
Ubx7wo2d5wUldgIiVot192WYF8BwCpGvUbmc+GmOGTeFzKQ4eMX/q4fxaCX6/lNsGIfo5jKId3k7
Tn2ibMD/lsyLX7gOZuw8daN2W1hTrRRb0NMuhT+ASoCXaCNaN2ziyzdg20ZuAlShl25DGbNM4NZQ
IeRsGMTsm6eWTl/GEDBUxmoDgSGT9LINq7bYOs5a3K9EluSCp1+BZCMn1xxEeUtEEzNibOlsZzfI
QsAaxsRj6GAawegtfQt6qbYn9GuS0K8hyMt/M8k2w3Ur+9JCC1w/lDz6r9gEd0poJm7pSN97sAfE
oc2Yuy8uJ4YyMxJLzoI8BHEjpJAp6JMkaSmtVsI6aEDsxU8lGEgCdPdggdbf1VPfdnlxIo1JBl2J
uResmlTLwg/lA9nRwrrL1aWDhbIPv9LHLdLnWZErjY7mJ+0B16M/K8AK2FPJSEfCovSQcKtymFJ9
kkV9t47DvLD8/YA77DDNICOicIY1fHEQa0YtDchpQKRRkF2Ka0+QUb1hh/IdD96uAPNWzL0eIYx5
lsIBDNN/7kqhOeEcs+BsK3cSgW4ion0WxFC2W1K1XSSdlsid/jcr79R2uAB6C6z1thlm4eNsZGRs
ImHhT101gvrjCOvJ1x9mYiMbGjUcIpr9grgNQM4ShGjZyGODDJ5EzMnM9iZKQW9ZHC8UQ3EN4fcY
JWmH/YQ7/fZihs5EWpDLAp8otZRyDgjXL5y55nApgM8toWQFKwi5MYMRsHg2XSExnrHqzTeoMcW8
VCKIsk4VBgO683ljjuSk8KuQ/uOQv2F7WG0qmYlaz550xUP9vO9InpUy0uaObuuhgE3lbXbCIEUf
AO6soVhlCHoCGHkVaMIn+74iLk0MNNuOZStj8VEMFq9Sdap4eBPeIsFuTRqo0VMSNJsYv6pUJBRT
99ax8ej+cLbvJ3iqKpH6YjUV76Qx3A/i5uUQMtJdHuqfyFF9kONbYWqcKgvjyt442vImAbrSWHIH
qY7hXoZi8hUtSeRyhCn9ro7xlvpRIbjeofO0Ah1TCy1uwsqGxoIa5Meo9BgGbqfrcxp0BKgsG8gI
Mwz8n/9SyFBDTINI7jR/v4TmVm0IGM9SGGqxk6FO6SjEfR9qFuAi2V2vxRAC6BJlR656+ml/8VqF
EScmA4HYWWcJCde11ZVkHutUwfDnkpNiA6t50Gvnf3nxXweRjUqkwL86iwliEfs9zTqFMJYwp53T
Iy7sqZ9YrZ1g6vO8gJEgOA5JyssTQkhw+bItL6THddZ4v1kmiGL9GkGVzCBbxjvtzyBnQbjwAGKr
/sgO1UkjwkRrySPBxeZi/2/Sg+oKYUNjyIgrVoQk+d9hEp30r69NWXZgPAVYNgPQo6OzeVtwrZAZ
bnWR9iqWwd2trRODj1iDq1hU8DYjbL4KeKB95Ex5XqErVOQ+EjvE+q6kVfaBHjYgvAmD/8bwfBKQ
xMTyB/iealTdlWGgqMkMppg6Gb03ZQT0gxuo4pfdMsjAfSD2bdCc4gCUXOZxmeYP5c2SlNGjaaje
YESNz6sAwft32V28M1iRp1KZ1uThn0QkcqYRghpMCrcp+OpCtLyv+DYczgB/V0aL43Atk6d29RAh
blSRD4NAsMBXCCAW+R7rtvFpy/zRmuQc+rWSo9UqC9r4L4PRx6IdyhLLwOEJRB8Iys/ofi/MebC0
tLdzWB4lbd6AHyf9IpxaTkGcsDHWXgBoHshPT8fJqXID57GDuQxIvMRE3iMpxnbkbEI4X0kIHOHi
GntA3ztGRwymzKTQMojyiLz5T5r3IqkKFi0jiYiLH7+NRdrQGakN585lm65E41PdSmny57eU/hvA
VQFIQIgiE0GzWjaIJkYbbs8MDzyOJOdDYpGX1TBV1c4KdX2jsxy9KTtrYDQFc/v6RxtwQJ8LtGCI
A707Uluh5MdYHoyFy0M/hiXmT9YUTQCv6MpzI8KUz0kfbmV/XkoFMy0iBshUD+nhypL0M8Pb1ZL7
33EVwIsrch8AhvSPbQj7beoadEfXAHbVsMTtXux7YFO7Ei+TwHh6PmINd5ptfaOfm9FBtDFGR1i0
RLsGA/BhrPbIcH/G6yIPRnXl2UMz5PY9vBF8UgyqcEVWMZGdefRv7bFciVo7J/xuG/H3LCTtVxdn
GMR7Ixiw010Je3xDAsk4i6YFgN+IYA8YrnwCD301ZMFSSR+vrMNwsuwebA80s5ZCaEDv4//KkuiU
CzJFot8R4y6YnJkFZe5mmcWegG3rElnajESahGL6Vr5SRnXQ3ilafWmHnLPOPFQe7wiV6GRrnuGN
vpWCcWTZJm0ZIyEu6ckDgnEOJSmIzn3/0m9M5WGWB22MJ1kFF9Vvw9F8/eag6BPSKTqTqEUcgUcI
eRLJoQK3PhGYMJ6rKxMJ2rTpDVF40v80Tjl4RH/NwOTEMb3kgFFuoE7BkT9NdmkxQr17wnqf2XkO
TTS643cfl5gS/IPpLbXSAfDZmTZaD40HUrsN4tP92V9igJaMBje3TUioerVV/H91tSmHjdeaXChD
r22BXdTQrKB84LF+Pwx3bhiCqeNC/8xG4jlrjm/MAdI7raRHMbBc0V6eqzUoKsfOoe5EtECz4Cka
gEF0yA+xzGWDbVniaJrCcMgWueVPJ31ny+OzyAetFbfAhqGUBgM9Zqnu4dRdpM2m7iZzm11QW2is
2LRb4rO0p7Ocw9EHlXEPVvxiQKDyRpyVhCFe5JhAVWTsuian642Or/h/jP0QxUb3lDgsOqeWllFi
3ULbIKnq+DD5qAVXZ7RTkwuKbOlG33ZBVVmrRhj4LMtM/2DjBPqghDVq4a5zp8JZwQDVmx+Jqvbp
0PsNzZuC5wqqj1BQ0FAqTbjH/H1DiozYd4cl2Y0TrAcBtd3bgXhFqVhQ6aFlw6ozhMcEzfcJaLFa
eUWta5DP4o9BAgd8CatirnmE8QDl4HpMdMLYVNIf/mLM6epEaKmttia+VhFYYC7i+q/wZf+oVVb2
JH1tzoi0OX2uTZKlmM/2Dvr7EPzR48bKiTNekt1/iXLlGM9K5rPRT5ROPaNllpT4v6Sectu40a7Q
X8/DjMHk7EEFF8aDPZcDrJXuwX0Cwsb9ddODINdhS4dlAvbJFO3kCDBqCCjtY3lfY0bSb1Kw42yu
jriveSiMgm9GOZV2RTCG01kgSsgQPjbPN8aLCnMurPuJZwm1lcPlHCsLTUraw1YuGu/3uZ8WSIu7
ZEA794CNLTSOtdmifWH99PMkWH27TvlaBz3shtfQnRZ/xemD5CT9Vujj6qoGftpIOrxI3S2iQ1Iq
Y5PIJ7keIRFgDjBUJZSpvDUo4oOQulSgx05wTKzM3OJ8iUsOzitJ+Mu5aSu1npYb7nsVwvgSHFDr
Sy3/2fjA6QEQsrQS2BX3W8F7Tzt45X8tQFrIUooo7JwbEtk8ebZzF9Ng6xZuRrjMufaKcWT8cyFQ
39d39oiOnhtuMXHA1JaXM0W66dkRiML1A8v3uW3APF1jelCQ67y1g9eVh9vyaiA1DxIv0CjD1jL5
ywxYFKBKtg/cd7xtm71vlVuRvQiyhFaUM9B78//yiSVvd35/B0c6K5w2JIhzNQjvrn09JxKhdTkU
+TiGtldBIQ9wPhcz/Rzpj8+jwAuRQMxqv8G3PQxWKWe8JYeMO6LzHOD5Nu9+sPHRDF8MnF0/a68V
AtONzhX1eTPb8h3xqNRJ7ZJguSuenmbN8PXgZcCaGjfvsWybumtVR3z3HpY2y9j+7/BkgeVyBnYC
zWzIs+UmAleD83SoP6EEUOkIeA6MxXRk0MyJn13Q8G7iRpBEHqzY5d25SRDLJTw9U77WbxugxFwj
XY6qVMSmBoYeFCLsXFyXXangNdanDJPZOgABZcIYeSSArPQJDBrFmhv0ca2FNLgCRvBYDzfUJXK5
CLlU/Pqk8+K2FaIS6/DrXYActdGCGZ8hCk0sjuWi0Ll77l8Q24bolgec8RnsCmt2STaBm7E02GWX
sv974Sj49VWlOKDcKZ83hwm38RD4q/uWB2a+qRwb6lAviNupY91oJ5HLm6IadAHTH6cjUbiPGqZf
aNidwtUwGVyKnSfqgVZ3WKdHHIYokddp5+B75towOOPYR1uypoMUu/KQlAYWGsnQEvB6jmkHe9x3
9wsES2YydcgJ7NjD2Hu3b/zU2veVAmsfvUot3sQXo//vrI9syEOnqthqnQYhAANCktYZFngenhwW
WvM/UJIgmBCGx5zSckyP8mSW97/oUcIbEKRD5vLa96pJj9hVhliKdKTYcT0j4cHrHHRyGgoNR6XV
+3QX8VkJLgJwhMrUiNFHqdHlP0gwMrs6DvfFw2FGz+Sx2akQmwcXbsSsOvLWl3GpiZVdZVeJG2/z
XNoHy5hKz187GD6vqs9HUeYv6DSCow0Tjv1+tRpIB/2C79qXpLNWo6jCJsjp0M478ulzfgPInKgR
cBMzpXtPrk+3aou2hDbrpV5genHostWP/mRpDuImdyccIl2o4nFCNVZsOk4jR28w3ZFKzok7Suta
umxOE4PgsNMjVowQYhZP4PydCU6RJax/JVnTOk6tsRa1Yvz/Fjg0Z1xEhn8rOtgrpfx8zaICXkBM
FAOHMbj4j6N7QbN71czzrgLhRLIneaw9dW+kRETalqXmZL4DBv1miXsEJfgQFVm56PQJPPFNMlDK
CrCcbwAs8CqaP3qks1h7nEi6p8qUgVDBug03zNjvfsmo2EeouxxGXIswueRnLx58MlN3O/iMJ+ci
Dkw9WaYhUKaCX8s7VchcwRCXtmM4JtFbYCumhVHqyNOMB68GMEWVUY30Q/n7flo7zeK156/6eunX
g5UcvyCtmuUi4g4TZFHpNPoAyRIIgt6bzJ0SCdTHUzIN0B6X+iXECe41apfndOqS3MSh1eEQ4CE0
jtNSIqDskzhmvMoki+JkJrpbb2+cK9vRqw5SybKsh/Pnr7aOtbPipayJnWyR3I7Pvr9QTLhAJzAf
SXPiwA6l+gYtLkxG8183XEnI+kT300wiOCIfkaa5kmtFPVvJSOJY91Hcsbi5CNmE63vvvD+2kcM4
IURh9n5Rvl35HaL22UMHMBOvRbC4elQXOArYozRBN2iIQ6cvvNGab2gOy9JoMpAXMGoCwPvX/XCS
Nsrv+QRz8hAAQ4gw7hInSWW11fVGbSa1H4Xrrhqrvh5aGb0EjIHt+Mrp1/P4nZ5wC95wt6HzlfKf
VfmgYnywCdezZWp9BSw8jZo0dsEQsmF/sMxtkZlHrSo61LcoTiD/AvyyFKHei653vAQWbrQkA74O
fhK+ek1L3vXDiQefbQylGk9wLkBj5PT9w/JDAU3bVP/ezdvyAPwFVHI9oan/SFms18cukENjm4PE
/KgbemG047SsuhrhP9u1YpiOnPkfS7W1j9FlmHUcQfXkVA5wmQau+LxdlkgYF8Ai/XvOP5X4cVlp
bfiCkw2uM1N5sdZQWwlBTZo52Qri0M35Z7bKFVcR5mTmh29yUEfuub6hOXy4RUdOcGbzCR6BcFXQ
8oT4dxuwYi47t3QWXTiUW5fBv9aqt4fkb0sLx7VEygKdnHn85pB/fIqkOrY1UuYv+qWGZw0UnvtW
MQ1Ip44RKJMc4rCn+KffIxFs5z/FDt7ErcsCnzUaDDOXIflogNFfo0LBQPTepaG4fRwCaw5Y0P/y
6Fznn+iOCTgdlIH5jCehZTuj96hiCJsNppNnId/iNi846PJD/ZXVETOqFnl/NXayPQ0NT0e38ed+
L3EphQ0aOFnhoRLm4ZPJ4j7/zEwJ/gtmha/xA9AjEzDdWkwVukrKCkraj3j2X4KqwBWeRcQCDdCG
nSmM4EpGDwyc5Bc3BNvufQC6rUSBQjVfP4+/C41Bg5GSMNCOmOu/oqHbh9MV8oyGSYMhjQyZS1eR
AAZyqVabklE/4vsQ2ZfQs+IcT/mj4UM4ww1K7uu9F60qK0kRS9lIYFaLjxe3keecJFQdOhE9qYNR
ATZfA+b+SDojZAsE4aUebBDb+IVhcknS8kWNQHZqDSBM5+3vmtR72QWc4WM4Efj8PWxr6ejWvIzB
4KZwqpcNue2hObEFI85/aoN0tOoTqRQf/lS3Ux9hSipWI0mukt5Ki+M8JTk0bjin6Yq1Kwo5/4cz
jJ81cO0qXIR1jAkl7cjaJ2zzPc6C2wrqKUamLh0MWKI4ZKx5p2I8/wN2HvvYeE+d/hNteUpkVhG3
bVxA3OZl9g/DdshSNVMi6GHeisC3pUF/NBna9aSKc0C6DUdnz7CU/gg0mNZ8EITCD2l4+DCpv/25
Ox56V90/1LbXz0kTKD97LLM55RSTPK1iQl9lTNLSI7TNVGOJeFBZFRkC/Ke8DGMxAUAaLFnp1/D0
hjelVX/DLMuiFxlo8TgygS4jCVEpITGWZy7HaoGSvgf8oeo9qV8Z4Tzp/q1bfrhKTiLDe/6V9/PB
BNk6UWgdQMl0AzW/eapG1ewQ5I678NOyucOZTqK+HA+0QSjExf3OOqJDsUrbMMlpA32SGvpEkr3i
kBVTuOSfXz05f0kpisqiaR1VvxR4Ibq620BlUXKn8MM6p/xXlWLjsnPKqDMw4AQDAQjlBgnSeBLp
hXeeMakBdXeuaosNbKOBW9u30r6bfxUK1Z6FcPfKRfnni4Nh1fTIkwaTLovxOiptKoa1vgX2gpS6
OE3JLL8JEgOdF8rjARaS2ljrcTfEgwcMlGvCFZ2qKHRg5gujp/jV0xXIt/PptLVCIq8ZVnpKtRbN
ycHKEvR9Cm+NJWtjwW/C2wqJTu2G9WEA10R1G0ftHq8p1q/02C5akHjTvpRwPDK+oeTIQW8I6XOi
nOsVsClMOdkwdncdb46vYD0hBZxqenEDLHWSd2vJpB3h/w6KucT9A8hW9rv+lEeA7nugcHOoVvNf
lSqDTzSXQIr4Dsaq5MxHJarqXpreVnFApmgALd16Fbu6KtFv1A6scH702FzM3rUNz6aM4SbnshlG
ISxTlLSHbQwDwnCEjjyVaHjNEwDYK02hGBS5iB6FreWmxPC30jMthMl7GqEvGC9azhiwiuI1pwaq
hzpZtt/1LxTV91CYZWSOUXqFNcONh4gLIyiFFkAdEhxYQFmfLxKafPS2dh5P+HJAntspj67Oh1/K
y/2JNf1kmn+/pJNlrKHZeGKN5SBjkv4l3+zYWGvT+IeTUMAxrTdUxhlZNjCIIaR/PTz9bkWruh1t
WwB2CwFDa5zhVobv0vlbUTrZM2aBhJtVKQYnyG5VGdZmVs0DoyC57+UdoHE09QMackqw4KUDZXzL
JDuAyx+cvyyoZQDRajO5brb2yIYjmB+RTE1PyLAu7z8BYMgY6O5QDHF60U9ZoKZwuwu/TVHbHCmF
w2gGCtAtSya8Sr6ka8HCt5+lsTE6TIb3ZEw9ZAyUC7FwcxnDlPzh93HgY61wpHQe097CyK+y7gL0
HXQjChoXLLD54qDzSmHURhbMlPsmGyLx1UU4izvRJN1Shoxaca/8dg4WF4hkmHz5vjnIffn/xx8/
6aNiMxKamSS+n+UFdQuPskRC+l07td8MDUxsHCjLQ/TtKiacsj43naZEg+sFC3N3H07oXRTBLmAd
b/3/4h6niI7D9yIzqPpa0gJLlbkAUOCBx1jhgPkvheW5npnujAX/anLNJ6MgpKA1TYcKJ1UfxiaK
lqBYjZBJLRkdDPnwMYH4caX+OW1YZfMaT7KznG55zmcaL1iwgajJCxIC0rqXu0cQxH1Wp4qkuefO
OtpbuvgcfzKlWkk2u5QdvV6KxhBpF5yQKM1B2/693SklBGOp7BRJG+82HXyGo7ujmktNr5f756sb
UtZxJGJ6qF0ZOZVdgLrdlnSAY0Km/QT0OMgFpYUf3jqltMCRoMkT7OClsaoikjAtzFODFIjG1/QG
nJ+2wTi3h/oqwYBVYYo4L01wGEIYh9DHSCyZtURnPnwYIQk8LpmunJW2B6BVbpmur8QZRA1Ynluu
rMlk26sVRtFfKFijsb100LCmCJXdjzkaTqf8SJpo1+A4M2hN48uCDvTUfJ4TjakcEf02S0EbIVxz
9qu9BIidjOuifdAlDBwgAxW3tHY0kFgSf3VpK2PFDX/HrfH8dyTRafdWctSEb4IchzA6Qx1Byeji
3+QA+wIy/iHb3yC3Pv5eeTF+YygDWoNnGvaB1FxFgGLJje7VVlN9n0W9XvvFTe0lfMY/x+aRuAbC
Iwd+qIQbvFEf4QgSj/PA4Uue/qxtM55ABYZZl0H79HkJwixhC5LtH9NvTNi7s6GGi41GRTmg9gU+
cRhG48VnWoz9Svf3xHCDHodHmOpzUw8rpwwSWR5e4rVxrYDA051niNmjMI8pk0jcQTyXlXhmSacf
JeB340OKlfiZqibKDp1kTkWdG3c6ctXkbBYq/ElEJj29DmA6+DOS9comlcFSq9zar+ymZAGlfnX5
PLj1u32XKBe6IlC2FRcGEuokWs6HWTqyxMV4uajeljy5SoJG1WuAAbp2dW7+4gFgeX/NV+1jpNT5
WPQFLNwth+aWJfNjvOX6WXlhbKtVlhZoWZ0ZLkHqJ79OPGvY5RkDMyQpn36AWBg5qt8Cz0mRwA3w
KhcoIlWHgnh3DosutQ7w0d1BtjEbaerTH72XXLFPAnbVjbozHSpR+3hpwkC3pzdHJ7ikaV52bnHv
Yxsk8iT7L/Untx9wzkQwv83UQU8OU7SvjyQSnKI3N1BiDd5vf3Sbb8CNn+NoQ7LhCJ6s3Omac1VF
ZcxvzMEoozeq38mhK3MtMSJWiSoCi5KVHAG2VfCQR+QFnRWBfuya3mZHWBY/l2bnZtY+UmlAPGda
yA+ftI1jDlRWINrUmsity70oWB74bhA+QCvJSJkbnM75b4cgAB7YQaKeJdQJ26+AvqhwLrTHpzZW
1IpLUNeCFYlB668uUCrogNiO+ADM9v0kA7Vg6DOKIPJcut3KvDkGDM42AbYXz+gcHPZQV9V1AHbG
nqN35Wr1x05+R86ZJyjjKXabk8HYhIGYZCltnYTnyOWF/NEkFws/NfQFAnmPeHqjdyVU2aPnNcKX
2tLdN/ntdyWWrcIuL/vMJA0Aq/yYGLHbwd9fwp7d7k2hdnAtpJ4IP0+2nnp4EBnpupq1486227gF
479aZldLTj4JHZAi6IB4X2VRrf3mZCz0Z+a/X2h0uqnpQPPHuJGpff3NbDQ2wIo2l7nBgD3XNFf8
uMzt3sEQMBHDFG+ddOZ6YYHI2XUMGiOsnGj+SA/VXWAv2i18sM+3x8I9kJIM06YZfoYCHs7Jmxl0
dIubM2nlRqc1NiBTBG2VywmcQfN9GPjToJhQcR6zP9bcXR+z0hVr2oDl8stfK8c6/CyyTZJjG0Dj
nM6Mjs3LeZ9TvI121yLTniXgE44yL+Tz132C/quoz26ptzxabm2pf2Wr4GMzShO8H88SalCyAXky
O2PDcEQ0bSte0zY6uF0rfT32Lumf7XvkoY/pmyinCV07fr7x/Ahnarqp32FFMaFXvtsNVKmsWxT1
jZPnNjewb6EMIdIXZn282oM+f+NbqnBWIjwcaJGWnq5vONLLAtoLm2zh1XcNmFIsBqRTvVEiqw33
3WVvuFteW+SIBQd8f6ckG7akPF8g2RxwBq4JmoqTT+NDGws5y7l/W6O9JhdaJ3L6TJuw8A1VC52N
EbMyJYn0EdAkfan2nw1Ar+Qqvat0FGahbn+sY9Xxq0+3NBxqcbFtLeIbz1VfyB9faONIWB7wBKrZ
N6N0XpCYW5Zt/jFF455Z5W+NoFrd2vJSenCsS8c4vij7DvNLeLZXeLwSkfP5JckPZkQEzS/Ou07y
Fp41BINcFlqbxMkiV9erSJohz3iMCoe1d2GxweC9VWzpwIPKnIOYRKQen59b+CAK+bFOZkiGNP7t
XBWAJtGl78zv/xIAqS2bo1Yo35yMcUUpWyUa1bL9CDCFaDmnXf3LJKJXfM77EGKQs8GLKxKrqhLq
c1nazMblb9waJWxN82/PjpGU5gHcctI3SPuexsM7Eu6JDC8afamoyyVrkzJV6F0n5oyCTH4uojB8
B0JHmq/lKVJiQoAY63N7te/ftW/CXRKW+REeF5eRdkcOyG5pmlcwUUITUiWG/SZJM+y2ufLAYtt2
dufKCgMDiVlFBYRpdnBJtKKkIq2qa1Ic6RCY0MxLZScMLt+MlyNFo7Xo56gNKZbAbk/TJ0VWi8mM
KymCkKSSXHuDLFJB/YNKhmo5z4QDpkR/i70v5REYfRG/1KmotpK0Daj6efaQnIsJhH4fy9g2JL34
lGvcx4CsG+xX9NV/trAB02uMd52WYO8tlKyRPQcTfYNQxa4XFd2LQkipgViz3rFnrfKIC60QHTSA
qcc2ih15sJNW98N8O0E0pGtBdMKBVmnDjyEALyZv9M9i6pyhnuT1LnjGLJBlMJpYJQxq8qJz85gI
57vpPP6NJoOXro3XvZqZ/+S5jrjkS3oVXvMws1dkmzz0AVKqcITeQqKps9WJFMY/1GeEZrwT/Kid
RhnoAWbLOdVpLCI1TMppj+cfoD/k+fDdPV4BsqAV9cSLMX1R16kr4k7TIMhbLycWhkaN4S/g7Uos
QbNSZG6ssXXJ2scuw+EHPIFt/UyqRIIJtYWf64UjKOzibtStrqkeZoELA6jwVeS3+enr93MYUmsQ
moQtxpQHY+LIH6IkuoiZ0DAED2CSB+vZDjHyEez9w4TwOhY4UTWR+5qTH/mSQk7VwkcZ+1Yy9TGi
cE8bXsfJGhrhzTjBdeHpV4hYspRNSa/ZxLwFkxQi04fzAtrzS3dHznMRdYpF9XphSEvetGs5S+0Y
bBF5U4aRvvlcGBo+JfrshniO9k/OoyyAP5PbEkXy7olLtwqpJcelNBmtLkqswbphWerpCqIQasRd
KkaCoTLWoKmZd0uK84Xybu1tQ0pYKnlZWv8GzRjpyD3wZa/2OFEh7bJpDDuyvKZTu7x2LIARAUQz
2kj29c3YcEz5fP9jV1E/86/79XQV2UbrUhWIfGEZQz4UaKxH6hxw2TMnlQr+8OGf9h49IhQ/VInb
1PUeg4ymPZDGVx0y0jDc3/XNJbdCb6DQcKQYZrUZhX5g8i2eaq7rzNX4J15hK6g76W8N3Ax/tWc9
H3yRmIIawCJxc60ShZ829TSn9IigURBk77dwMQa2Ed7INE9xRI0cCdK86q6BXIO3yPLVEno76D/h
x+5O0gjG3nqS6UOMkuvtoswk6IDEkbVMQbQxPGndlNyBM+i+0UhIT1tldbLWPQk8d5Scl7yWcRES
J2RWuLAwDZN7AVrFCfrl9hkGk5Xz3mlY+qefgriTeG/u9IbmT5zkzJv1cs6GAMGawr1vKt+JA72Q
SUDz/IvJzOyuv7+OqideXlCxHZ/QdtvzXdqe7skYRiT/cOZPHiy4goCgR7qbUALhyhbTz6YBmj+1
WaYZJmAOSSG5rlDalo0QfXymfb71hMshtF8BKzBGDSYryp38QOc8Y2mmPdATBYa5vFrn08oljvgM
XhqsJMxALtRv+pPID4WyEbc3KSgJNpZg5WPfCBA2+whkHo68KBwVwT4+0V0ZJpKsEcXn+rXS9Ihp
xDq+P0BhC4GaSXlkgtM5nyzqvzAtM3uXBtVQZ0/Jum3XS+TcRDkTlQkiFteq2KT0GP4Ww0cbxdQ8
cVryllHcUxdXG+NaVPs+WYcX0IW3qaf4J680tATxznK1D4KxQv3yJikZsvSjohlAZ7F7d3H+YjS+
EM8yNUf3yDys0GUEQYuxLcyGmZBZFkbbHWIPlaq7N7FOP/gdcW77NcmArofL724HCKO64txEmLiF
ivLqwauPBf87CLPWTfwuFgwydSE0GrSsPLAUsjhfFJZ5UkpkhhckW8c8jPKMbjAEExR8BU7K5jmQ
Yn92ovnD2sJ1rLrP8nPTq2IauIO6DDCjhgouVppVXTzqGItRhyEZD4Ag5hUbZWGFTJW2xs/iQm6m
rktLX12Wqsyhrtd/tz0lPS1Y2x+L0cXi3mS8Co7Ecgx3UnRBy2MoI2slGWxzYOavMqcbzsRacDf/
DOH7lL5fbaZ1eDHpp0zsq+uDAQNlL3FWKQVxaBbJbMF7n2mDqxLeojNDN7z8j8njeFUm+xx5D0yw
m9PFvykNHsuueIGWgce6TlkcNLj7BK0+BNjWZNLNFFbGZyypcNJwX0mJHdpPuxI9O0FnCFYhgSCn
X5aWEHPumala7kBBswn6gXrQGjEzb7PFK9W65suBVQzd9QMADgG+GNVF7F+B6zqo3TISINt5s2oT
igwJbSL6oRqIp+kAJKmIUNCeWNIU3xPub0PRp+eVoaSSpBL/7zHTGzmXV3+RIM88y8pjUUqXRk6p
qQeqt2FfgOMpif+Z42CowTCMtpnu8XD1sbYHUyOJ24p8PHM5LVMcnKyDwoXG74sxShiU1tptxgRE
mYY1t+N1wGpahrHXxLxlS9LNMOHLPA/J7CPf3COlogYY72bqYY0io4+jE3H+3sw5Z8IdbSU4vAKc
6VBXVPUmrFD+pl7Wt1GimJzmxd/vU1T9qXPo2sXnbwK9Zhf2Y+Gp/miJSNv6kSBfgA+4eSIeu/+L
630sDciDnOCjvpgLrR8Y59NLpS85yE+3bSI40nPj0UiEus5+O7pcTakF0IQJEhoY66+450+qtogc
FtHudGGiBQQcygLYGEX0NTiWZ+pF6l75kxPDaA08QhOsb6zS3RLcB2iZ+/ol1GIIp1wbHpktJyB6
wdtjUPAk92JU+AkPVYVCtERDpg+4bWW0+0t1n323uFL7jV1PaXL10rbX687YHKMzgECBW+ykV0ep
VMWRXPfi4MhVEujrjzsprQ+TAWwl9r5hNYBh3osynfCSAcY6tCP3Hn4kBz17zkeskj7ZysUAHnoK
MpypYomZxlI66GCjZBIt5JLAScfgeJ51PpbrLhwHtyVSZvFN2NGneToJY3GsK57pe8/F2Ro1Ww7w
VGiw7gQhBbVNbVV0k0+scWpPjtZW7aSKC9L1KuRJ4pQLx8qUZFIwvzoFO7gTIKMmhwedZQzE1nZr
53TxKQkFgLhaclT4pJAlmnZEm37c27APM2LoDNaDZ2wCUfdZrjK8jGcYf+Sg/HQUGFoNzHrQJRv/
aGEo6wm+UrEDnwWXkI6+9yV+/1l9u3K2dqxu7eTvUkVeGm3K50r/YQfQ1h61Oim/dm+S8FEM+KuN
qiMHHlK6+940qwCRn4+8KMqInhArgHgiw+fFZb71iqXJ45qJYZYjD3m6NL1HdgcNLADhYxZ89ucO
SLh8ZhC69zDndZFPpECkyj9Ppk9bzZJp70neZw61og5PhczhCaNjUw/PsO2jnk+HdUTdZNapqL/e
W+W+2NQii7fmxnwepgNgEgcmuEvCy57ayhGcRoMUTI02TgJJwMik3oMHzuB/tKQ3cEE54jXt3bQc
RgJkDMxD1jonYQ0g2VVufpBt/Uhp3OrZtnl+QlChu40K8r7RtjAyGmChsq8yVYhZvhEYGxfUwVyV
rW1op8kspDFu754qKkoL/K3QOjCeiQN0YMPPJI2ohSHA9WTdnaanrbJBBLaNEioqzyMTIdsDT6v1
9Ke8WwpLvTxaDADb0kN4rfBbOTAw19XeJR6G9eBqQd00a9BU1zWN0Q/G9GRx4YupWEunGDH2S4MQ
uQJhkymzadQ+kXPLpP9zScso72ZNfy2UDCI0dR19GzPI+wXKg2EufdGTiwmz0xADOgz5qyoZhQD+
65W5qtkdltK/r17drkRPWBekXX9PUgpLB8lZjdNBEIO8QKxGPObo30RcVFkCTCO48Kj+tSvMld5a
w6PfjHRO9cQvUBsgo/TMRG2QZ1A0jCUf0lvKed3ob1Ybm51KIf3ySdJrox382kAf+AusBIqPjos3
a/ZanhIOh4IUbE5ivp605I3s3z7coRQvrxd/6azfXCXGrT3XEj9L/n6og4qtW5GVW3bFwwfQvKvr
FjKabiwnErPvZTgzrm5swRGDqi7ERQMg6UJSCRFv+w5QlLa4umkdz+KTgsgp518r5AaHDT4aXL5z
wJdLpRwxNjovac291V6h4PGNj2qmHRGVPeDWq19R/lj4wqTnJ56Fi/59Fuao72w/C6PvgFijep2G
0BFokgiwamzIJVBcH/9keIyTMcgQQNRjlfPFa8dAwgAyl8x3ahDWP46+K0nDy0D5BnFzlew0AyiY
b07QSKWNGLpX3oe8kk5BXhnMxlPzhExfRvJmQIfkR5ADts0XtYEY9+n6seWBE7OufIgIbU4IN5YX
gh5gDRJ1lrkKnIS9Ccq8GBuATRlE1ha4vf93vGgKkhkyUCnhV/Z4vVkK4zNS8lMuiw/P0dWBkwaI
6gGhP7ogJBaVjOtDrMev8/Da0m9Ca64eX8vtBEnJw+TefcSnxujWSTsWdl8ChTtxrYV89uzi2Rc1
eleemlJ9rVb8hjWHdAGH437HFSawGR946aVCu1kbCuG7zhGKy7kryhoRC5+g5Ph973RP14IWCQBF
jImchTfyHHkigM0RRIfsAWiTAHcNjdGNcZOhVAvHNuq0n+4ssPnhNv/u+KigLToFlGhmJ0ADFU2j
FZ8POCVk9PTA6wDoyGxHsM6VeVMUn+40qp8kQbxjajEEwQtAulBXyes7W43MwshymUqYnZn4ldUI
27bxEBzRrveRbwZ3h/YtApVfswJFzGqz9pUAESqwQo9zv2l0aMGhrn+n/KJyJyZfM3gC8BqFNH0e
mDvdwin4FBpaj1lNSKPDnqTv/YDIHjXRWGlz7zOq0V70TZkgLwrVEuHES+WUeRkf6FD3MadNkpFO
YuMJw0dKeGZ0kMpsaGY7evV5f7/jslZ/dg9TFRnqY1YJMmTgvCGfNVpM3lQyZ46jhK+QhMQmfoTZ
3yXE0SBzkzG9mEcRKEuI/ZBsHft4WNRBIEJcVY0mEFYNgbJKSiLBo185gZLW3+V0D0wjYBgPFvmb
U2GWMrL8VmSQoVJ+jVtPq6kqgeIIYWFV504jh53DfRo8mFY9WtMrKNvUxle6iLoE64VRyPJyRGOu
TS4XsFWOkIvswal1RYZdC/8vdJ/QzJF92lBRPxslj/OKNEHPDc/G3IQgxmvmglMBPVCF94uS3Whq
cDLq653yI4wF+1j1z/StX78PXCSz++VXKnNbKS2brK2I2boFMtD8sD0f+Bd2ha4Eh15kvTPK73/a
eBXEoJkO+s69/bfJJR1kh0nH/Ky85xLONhdGzZTohz3/B14qPJrKre2EPWFDNlZwldNDziBGhJVA
MpAZcpXNZGpdClcbVCcX49rP5ZUIhNL3Y61v83GGhZ2m4GTsj8yJPjyRNHjoyUZpuo0e05KCV08z
1LMelBFdDIC/bb6aZ6e2O/RP3Y/9YdEMJGQmqWFSjGrsZabx315pbUJyx+Bdvx9hAUjRzDcayFwH
lugeJmce7Z5E6aIaC07UQJecePLe2zBicgR5W3myKLgdGP4PDcPMKGGMoloOADDIjc6+0b3l/T4T
Sdix/ae3H1g0k6x9LcEzmOyBilbkguqKGDyCWKyBryMl7U6MdLPgmrhpw/nSk865gwuRQwbIU4Ep
ARSqxBrqkAE+QxMA4O13yz7iOXAEf9oVkqYgxx9IrfbpbxjoTTPZkQ3ArQ3mcPl3vrkBcOmd6R03
8VL3AAvXoRkB8vMpunAZlWjEzCnkfgEdmzwPXG88NWC/BGc6azRm6NkYMR0IBf+cTzmUXxWjVl0K
jbmwKAb+JGyw2LmFTpuFPsBaQehA/7SI8ZYj3kyIWrrKqcrRHuH5Of10CrpU59EIrwrcpj6Pm+Yw
GoUk2oTbfllK7Ao9ycpE/sf5p3Sfg3XXFgCpJwdXfLC7Wzx0RradMyWvcHv20xOSXQWpefyezkQh
CanoOiaOtsUDRjSCfaEB+2SD0k82wnc6HC8IxC8L5AJR8Mkt3oHDTFyeRP9OmDSHnSZGnrFC7d88
4YgbErwXijvBzIkatATZJq/hoz+cEu9jgHXZnMKrLdqG/gJVlLlkzSIQuPDTfl73qYBDK3C0lEpq
SNylgi4WaK/pRctk8DyMEiJeVgN3PqxU/t8CVml5/BZlPaG/FS5jX3hag6NKqyYehz/dR7Qm/OsZ
td8eh+eDlDerNHdtH5HxvQPhNS7JlnxrVuNCCK+ABzGx6bvgfc4WqsXvRfGnBrx7Jn7jeJV4ANnr
MPHvH7hne6iZms8PPbHaJLRBL8VWhmPjsJHBpyYAzK6mzKQrtiAfa4wWAfjbVpyl4tn2JppE0xBp
q4+BN8LVd7V6J3fG/lXPMkCzvvfvmLi6CJ77IicACvx0S0DVpfArc4ynAj6vms3wJZHm8I5PgkQ3
meNhTCk+OhfUHJl+IbkbzL0JTCjiEnPuvqc708LhG7cHk63mc5d2Z0LMmotIUKHvZyUnQlvuhqyv
W26tag3dVpss2XhcL2C0pOSJlWWJkDx2kmBvYqBAkSKM/V4dGmPYZEcdwj77CVBMxCylzz6FD1iE
jXUvFgmnot0lRo2Lg7Vdou8aZoR+OtintQ8OyHfZ7dBOxg2VTz8lCmoihaGHo5KiqFyhO1MhQuZY
nJes7sIUCPIDnLq0lM+0nsrmwc3xafVFwdZGAG0x/sz3SHkTn4pHmiouXfFV+X6XhejKCxkvvIM4
QcFOloVY4TG3/VG+IAO84n0flU3TOHx8qayv9IyrgEl751O5MGONqYrn2P1IoSRXV6f9G1NUekZx
EnbM4sFIqrF3MGx6WCTE+lhX+LVPaC/hrXe665NqVJf2fTi/AdIQ14Vj2S56VjtvvsT84P6cLsqI
FH5QIajXbh43B3l1ptdp4fSF1E4mU4FZEAwzSeXCTaMPCeNQlJSjSJHFaXTySIJsGNHIMd9ikliq
lKrMmpAEtLsnLAn4rxFEL7zq5J8sXzWqVPpkBOBJQVTGL1/u6V7CM79xyU4IE3EFnHZe3SmUQNyO
ENVSEQo3ODQTQyP6AECOXZ1xV/lXQDhxzGOVL3tF2FovU8ULN8dfOqlhDyk74IOHDGYRw008WBjB
fCCkN+xXUV45+9OjP8CujiOD9C2782610pjTYt7X8azHFwK8CMggvJ7DN/C6923WLQ8V8wmJOETd
AAMW2tmImAkU13OGdnovBjCfLiUyfQQQoLhw3QVka4P6kcdwi6dmK3TICZYtnVtJb6Cfa8+CbKS9
vpzfC4SZrjlodVp5DPcNl+1N4t+qHBjHwegPPK7IzjMOQauWVJm52hHp4Pa2UH2/hP70NRfpXNqs
AIu3wik8Pge/eo5dvbiuKoNGu0QHmNVWYE8jNq1COEsjLk8GdxZJlrsEk8vo0iYu0mBR/jvGX8Az
p4nFy71jQUGD7LyQY6YF78L2Nq7Hpd4FL6J+hRVsYEf0RCa+5zt1VcEhc6MSrM5kuuQQVnzdOA8a
1gUTkOQNe4M6SmwbPIQmB2ACThWAVYyXaeznEQwAERZZ6eQd+7tsHxCnSjfKhwIAdLnS+OmasGnj
Pwcc8Rl3KYzxTHHnisXOOFtAhMCnU/KL7FycdOm+wkpzmkCO6Ch1U9/nPZg0TRJHhIRaQ4lG8q/c
lXYwxy/bAUwyV4WhahnKabBe2nrloafbmX3AmXjlu+UWtQ2tHEOFBkNMJ9IXX8aWI+W+CfA3N4hK
4eqozxkuaJGLB7lga9zA6EBs9XZi8c+DVV6goCq9wh/tceNOGkaC1hFRScbsy6cpJ1qwe9VBhm79
2skeYPkyFGuVHLoCZ8TtiNFTiu2pq1f1sUIvYP0sivk8v3fLw28WK0ALpx3EY6ReBpHq27n0FD6G
GVT/WcX8bti1vXsAXNQWWrl6WFHn3JiuFa3WYUbLC9ooHZlPe7r8784TOV/Ft3sqQhqgiHV+glM7
sVbAuUfhZn54Du4Eq5ktejFSvMrcBZWmBGMLAFjUJkz/ylwXS7u1PISffmEQnAKkiScMQhKsCX+N
yrmS3f3W+b2nRecyrdqus8xQts0SM9Dbc4haaHHkc8nFI+uvbdwunHGhhR2o72NYVyIprojeVdYa
R8LN7fAZVCdC/Eet2OMtsnqrV9h0P8NN/TKM7tM88hZXoNuEP+YZ4jFnrX/MblygpH1C7r6jvoHH
VELN8m75My/G0i7EGgDnBVsJS5+OvBc0cpBz0Gk9CignbtiXBCwRrrR2L2yDoym22uj7OLcvPdkE
d0L+VP1wK4zHhU5uFLGhMHRDrdLOclglCUzLjvrTEOIwG5RQk/hUk+ZECdiKSkdizDXIaXkKM2gs
6ClnH1unW80TX1x0oT2kG8GfbP5ygJoYKBmd6eozs6tOxJUCHy4Fv76WjGbGC2jaVECMfy1n4FJ/
lfTkws/hdOHmKOhXjgnati120weROn99pdRJkWSGPltHLPc0bTWitHcSifcnzIO8UziQKoSS5tVN
9YWaEFVlVjnPE3HX75Rbl3LJBJs++Pwi652Lvw9WUugwYaQBh7ELh1Lo7/WZFu7lB5qy1fZ1cNUn
S974NMBe5HO1d4veSfDRl62EzA5KQspMdjtK541fs4/OaUrZjR4HJlg5Tg1tEoHZsXhOayujPE+2
DDtaQ9WjazzdAsn2sYMO5h8YpMTn3S90qJY9JY+FMpYBoaZ/qukW6EUgfutLU0t77cQuUb1vsOz8
mzeDrCFeBBm4NpZ1YCydGh7fVoPP9QoBDLEcj6Uiq027LO5ZjgF2zfR83zj7yec5bxFh9xyXsv/h
6BUkNJFgXMjKCshrcMaa3OL0lrA/vsRscFQ2K0EELjrApULGFJ4rRa+r6EV+Obh+oE+iPOigIvNm
Ox01Dba+2us2fxFfOxmdnMiaivuEHM6eHrPfbF23HnW+tCz7/Q1WCp36/h8hpRxulg51hnUobDg4
Ye5y3b0w1WpUCbCoKUflgmA3Kmg3HeqUcTqGQywDNwUgfUquyTlijGs3J4BMWMXsltJ/VRRQ/rpr
03vkWOUXP1kFtRyEAXgBS61c2vJdNYCbgtW8AxIW3PNx9VUKoOf8XTBcW/1FfJj8mZ02yPMWL4Vw
AUX6Bu3O1MrYRUxeb6/Z8QE5XUdgKLLMAjOu5MKP9ciHfqSPR2QpTXMmqUx7L4eJtS5n2DtBQuAf
K91KaIcnkqbsJ+go+9mzFRep2u0mJYTmC9HNHrfiKnDhrDA+J1uatCnEOgN5Awyd394+D7B2JVf1
kffzAPEJ/3oM6rFWuqS1nxbnBMlslc4KiWxG/4rQZZCV/eOP/Iq8BS/EmJHc0cK4Hpg3YnPmW7Nk
FbgjZt/nOWjzG5gI+bZXWFSKJOTVqpIKMTq8DhHG2CzA/8Opy85lyDFtTWabACHvz8w82FUT2w8O
LiV2+YC2n/cXBm+8TDlhYBYKlUnfu/II1uvdtAYoTQ3Hwq2oq0HvZrbxmi173Ca1UGyVaFkhylRU
yYO6Tq0qU1ztTrq95X9jtHmkS0MueQcBRN6rSQB2/dkPft1FUTi3L+lRAsVpH7riC/uySJ5cBcAG
IcON4tYO3Hs5/VZIg+Ut8ePJUJDylCmR6ssZB/ymNccjLKYM8KoG9NsWJFojx6tVAjCpNjx5ga54
IGOxdecBzmKC+cMS6LF2o2Hj0tFqZVQCyOwd07w9jn89pGG5pnqqqVjRjy1aE/T7zchjwsRW04sU
077ykoj6Xw5ijS6TJY75yh2jhVMicNoAjH79v/sjCyy1pIXvvPxa1hOqzW8c1Qv0/3W72VuQ1lFv
KuYICE0IshVsl2jIWEkt/9zl3igiPLhmsrV1x02jD+NjmbxNiXVGkUUv0xlFA6ps7zZHMa+t76yD
OqPzLN/5bl2AzBKhSJQTiodLLcKNONfpKBqIZebHzIdQv4SehTcRuUXs1bw8zKms6HUt5KDSWkhR
Pf35fy4Z1Y2nm2twvdeZNzQa5HfMCkXOoHrc5K5s/FQdUCMwRtsRvOhCDcHXlodHxB5FzRRAt0KS
NmkVyGamyEzAR0dai5eFc8vkYGCNtjnRe8ZwSw6RJCFm9EZr1GsQE1lWvXbHxCPMHYere94FaR9b
njY9sIqhOc5Rumbdprp7lL/uvrrqfj9kNXMWfEIMx++TqgzKD96hMEDkxhAsZFgbqyYLPE6uOZen
YgnonNjUhnDlJ5HqjQcky52RcbOI4fNX0igT0KlSTml7H6uTY+rbP6ydwniewNRyAvq2itMKBhf+
er0qGaD8+uy/KG1ljrMQaKxP7rHPXQOgY0SoFN9NC0DR7VZGvCmx2jRugN25j32SXEzW1TDpv1Q8
6XHUfHH7pv1Y3KTdxGIM75wBzpa+dZGPDERMhkCf14JHU7oAtfvF3r1nuJzh0mRdNR4wr/fCf92B
A4iMbST2gdesfd03nm0oy5XKvngqvdXs6nTUbklWu8WxYvuPwUOEF29qyXUxZI1bI5b4HJaLveYl
LOHgmLT6LIiX9/GwrbyR5uknwG9zfCYrQ7oLKHwepx2EY1NNSQ7zOIxyzcRpV6xOFvoxXa/1myWQ
EdQqUnEwoLjjAGvE6J4JWZSitJZ8Lx2fCvtW4PusDahgVdWM0yszRxtjTTaWmyYQDoeIa8VCdWX4
Jsx8wrlMANoljXX5zE545Zb8w4EgbKHeIN8LMBzK1zBiseuHijKcBn6T+uyCdvVLrLMUiUUofoQ6
wTx1bEOejh9fZj8tzyuPlhtSWa7JjhUht8nMZhKWq/higZiAdU3vkz7I+34Z7MPNZUrqdBwaB9bt
fyGYLFds6Cl25coO306gmHVA06M8Xvw/EGmY+Ran1oTRJoCoVzr4B5kqh8zzv/6Y5DfLUsgA+kDa
HyiBOMkj/muw6KUH1A6OrlF1lDnc1++h1CIuIjJCINaJBG3Rp+ez3DSQbBcz+2kJTlCRvobT1yc4
DGrEgDhgFA5trbo1qhZcEeKWoJVhd7GBv3RaVUKsOhl7I34RRu/obqWztBVAU4rak+9M60NtiIv5
K7YR1cNMBHcEQgJOFMcSaVCXxmfJm2Bnf55ReEOE5eNL8JpT4Uz/roKNVJaYKYSeLfg9iSE3qZ8c
0wTZoNST+unAwz4rSFHhfYUuNQfghCv8GNaLEAFWmZKlNZ5vWhbp4+sT0yO/NmiZxuR8revzgleg
4GcJ9XqO+kAsquQT78YUpqaWJ0Y+TNnHPrGPWxOYfQD0ZPB2R+wtSzat1aX8SYaLkUkvfVcvRMiE
+tVN2sd55NfqDeoOLWkQwwIc6+WGm0GW4UEwQnoYXpoKXAIT4xmnLwqIqrzRcRc86jtSleXCmRFc
jjygpyAppxDsFu2jgs2aFoGwZ+RjJ5aoGlRcoM2UxCDqlwXmo4daKTHwgE+vK0Bxm8OJSDC0yDFV
THE7jd3lwj6EcvFohr2FycVukvYuKIN/DPX5eg5x8Tc96ktEtuXFra3YkxIeUEAatiRElUKKlCIv
ch5UapdxB/PvG7gLChyF6bgnIONrLNyqKfo+mN+xuT2hHg1VB1+ITES3e5MSP7g3TWh4nBxG+Fxj
b3h73onQgQ3kxf6m1Uz/Gz6oyzAtMVyniP+viGiUZqO2/vwiAfwHQne63Rp3FcT4DcceweDKySfC
/f4Rfwra4ia9VTnt5escuIFG9dCuW2p8n0QLJRX0oFC+YtV7lSETCDpMdXJsZ2wqOHar4tWwjHQH
S8jeLwlfalgaxjVA0UCyXbK4+sJqwp28txov32yk6buHE/cvT9Pdg8T+/w6of3xohYMjBrH5gGbp
Wh6nFSrBeEhOOQ8fNhv9oSE0eM0MIEBTNblSGowhCXIC8+kaPiwlzaV4L86S8ncIuEwUo43sgdSL
6AltnJDsDjK0SEHu+K4vHz4q64AdqWwS2b0Pv9esM+6x+XBVvJ4pOG/iAat/XWaRBPC34NlTIH87
GV1s0xrsMofF/D6my8jeSNDxFpooM4mNxKg057QU6azdE/HLy1cU1zzSm5Ws4gVaVf+ZFhnHKfGU
nhOfweCeVsbIfABaL6sQWZVPIVw1k2hL+hAxFK8qoFFrQgQ2eoaT6mkPRfJyFlOR2PkQtoRlQDw+
7ivDAEQKs/G/69q8h8A+cdt+UItFEXg0kDUjDkPo94OnPxA9YQMq0kZDJEaxb3bH9v3p4WSHF9sO
qyl/fZh2asLw3rzNZm1/QcmpOSdiI2ckgfsYUKTN3M0g15ncfLmehp8ZaEFkGDaPyyVU26JYL8GW
HvfcHJxdWf+UIa/W0m1drstJALKWqW/MI87oHYGLWQOUD2EuJa5Ey3otAtT+C+HI4s8i/JIcLBkS
aFiTBUJaPmnxJyLjJay5fUUU16FQwKn8sNLZjD6OXcx/zqUDhp3jDo+ajimgm0zTWUZRnOcRMvoB
UI6JaZyl1LqVe8ZUP/qMVD2Z+KTU4aK0tpsw/zDWzx5N7pVBwcdUTlSxahQ4tB7tpctFQW/aAXQF
209snfSq6IIYtJwzG2F67sOD9btWqrtyNFDuvbUgj/FEF064EWg9u6zV1f2+bfK/KvP/4c6G6MJI
6oahW9+jhYap8In7gPrWzuuHxAmH6D5agSkIrrO+jBWWcksXeZS3Yc0wGWqEHZ4SyLrxI5DkER1s
1U5hy0rlCjmvIV0smnFSMYmkJhmLSIkWgOQWRK9R2arNSGbks46m1YHzCunyLA8bpH//qjEHqiOM
dv8O8s1CRWIaWXfYEHYPX9t186v+tL3q6Q6+E5sxMflyUX2oO4sZdG/ZhR9FpH0xzJXmo8Uuttlt
iNR93tPaZhAFxlGFezdzvKxlVYQhyNMwXGI990ZrKtVu1o2Wn+GrpI23//0UwYMETrFR0VqZ9hfO
4u0fD3YSykqCKiNQCbQR2RhzXiPhvdZL+LM2S+SpkpCr15zJxPi7YJXI/qS6T4aZIWZsOdH85pcg
Lmr+QgIlg5wt5yi0WP7fPtfBLKMZttX+xo7AqqkxZOQKy+s0ADlVazrseox7cmzZDqG1qIGKG6Us
E34eVLNlaYJbj9qtHVhd9UBc9S70M/I/GF5fJ8wVVxjUmPiamviUNm5kYPivfYnjKpQ9E3kcSx4V
vkRG1OO9NNwZP/nG3csDDDOKW5FpGl7g2wjxIrjP3rgTG54DeRloq/Be1wVfHjDO0LMdt6LCUEa8
K3O57e3tHZ5MjmZgJ9cUbazmoriuPXnavZVRZR3WLKoGx9GMhaCxxPrD1ScXSjZOGFzLOkQEcbV5
ZlYKssPaVVzDxG8tTK99ZcizY81FPdr7/EJnQLfyAhjIWKF/Zn+g/qveD82xOpmPtGEj9BX8I2Oc
5dGqZDWVZf8H+nPpOrtccHWhMiMruojbZGhyM1PM6dG7Wa+jsqUghbIWxlmnAS/IvPrKQbLkUiKp
q/lL8HetaceePIvn5nQ1PSIbUmtKfmzauvEwkgpCRh/fQrsqnV6/kVWkhBpDFQJkCa6Fp9GjKY2g
Jy8q34J02ftoZd2GoKvH5gCXS9KuV7Es9Wp8vCPufv9NvqkDi5TCPUr0a7RrWX6JXcQ1xS1ZyPmL
5zYYFStLv9sPcZSj7b2MI1ELzvD8KIvWNgmhAkGt2NeCxtGbAksR81fCNXjd+QeGv0KDW2e82t6n
OFHfuvix2Ii8cHQY4S2gfGH7h90P2/RHTYZKqFmdBKUuehWNDgmA3uRe8s5t4BGZL56SWr6OZqrv
yv31Q7rWifGaBjo67Pa8WlvDEXtfYpKeGImkbjXNTk5WGmyWopvPU/Gv43hMkfwFIy4dlbw41NFI
pfW0QTGftmktEUfJfGAwhHo3F9WH6vpfoAgslGjX125dWhcyzMODejfNpWr7Ria6UtNy/p2Sp7GD
bSgZwTNGFwdwNXnYX8T73FxhwsyZ3/CycxU3pV1nsHzaj3eU4xLRmXIk6df5ePs0w+7XivZ+HBc5
1oJoYB6RZxvA31xY/VGzfa/SmKcgl4V/jXwsngpD7TJReAqHwtwM21TRrDNZJNCdcHRhWUBuIt27
lHbKsp349UZMiPHJAlA23KjTQMTsgxMV4VTxSdznZ3viV72ced1cKF7Lusacmk8OgohDmB8iuE0E
ao5Lkm4I1NFf9nCC0Jy+HIs/AO2Soxio3+3DrGTXTP4I/D0jI1c4skyyMwF30z+ronv0tYELozw5
9Jtg3eu4RE3oU3+QCh7Y42+YfrDyRCrBw2URIkErTH7+oPBOWAllJdp+DEUwWAbEEPsbcaGfWfVz
91ZhYgWMzm0n20OERejlI2rMcxYDNDAESh9R/qvEb21C5kAjTJM0shnjPT5AWAE56jEwGR+ufnQK
JI4WtI4d/ifIeU7jcKWDAOl7/DPJwLFrQ/FHw9CZLnHsrp1sWBvfkYDUWCIzKrt9TrQTvzSgm+Zh
woq4ImjbWFj0ZpEgQ6tX7gjGkDZyPaeBin9Eig5jns/VFHhJclIc8PqU9mNc3LSDTaL99D73a3qp
R8PzldpJzs3YReTv6r2kLU+xsuYt4ciGOoCHPDKQCPjDNZpnQobDYIKi71eV+so8HlOWNFo5cm8w
ZpqbO7eILHtMlH43l7LW2WILrPZUOPqgIOCv+Wwt2uLDdJH4JdGMAE9h3qZ+SnxzF2rxX32+eEej
gY3p8O7S/XYaLqSqCfw+5raK0e0cH8mv5dCPlm2eXiBo5S3l7q8dw1zkaGguTR+62S6TH4XPYOQF
WDAEDgY2BJ6aa9yPgfu8EVvyFs5KlEcQvQs2v+HljYc5PfWsY9WKXMy2WiLgZSIjNmN9yJfYIfI1
CjhXiJQZrsBrh1JReXxna+SuST6XJXBATGj1hl/coKGfCRfocbBYYuR3WXb44XTv8tzdlhh0MZR+
GYTdZ2T8AO3KCIqZ1bLGntTNM8SQ+HyzIV00ftvZ6spmXRb1QHPRoELXysEknDL4sv1xS23Mf8U4
fn/squaOnQ5pabeuiceq69bPZBll/zDFxEO8j0YS+OIGSjbdspMf/L57TnbKYqjuUCIP5GniJsaX
2hijCCJcUFkqPPNThbV2WFS7fAolssWjXdCwKNYwy/0m+6BX84o3j9y+L1bqSjccoC578oDZQ7BD
mYVExPB8+fnC97m+ZkvRA1AKkChrqXMsFZPGZaPF77Bfb3nSYdFepEGbzu/MtfETQhw0AHR9lAcy
eB9RdJf3mLl5Zo5Lvx4Nm+6EhJiAC61xgPTDQ76sO6V66TxfA5iUbfBaRguxsR97DmHdeT8lQTn8
iAANLhnrzSiJuCk8Yoe7TTD8Q2CcjHhgPZ99w4nP/g7oXOYXGy5D7KFleXr18gvljtOc8Wucg0oD
Yurxr4GbtOC0XiFfTNdV9887hw/8IMSXuo0shkRs5c5TuyRnTtJ5C8DZ8yzNEyKrP3hCBHF6IJj1
eRcYtSCZDfbJfXjJu7v7mVAO0/QMsxRY5gWWG9wfsCdwxWDuqakYdBbB37oLVxIYpTTReSyV3VBZ
23jPW6QQXSr86CRQ50ki9DcFJA7OCpfFCcSfXKbHf7f/vziWJoMJcVq4TWcbqSLB/v/2OLBYrq2w
wAUfjWF7GJm25fI810Ev2ZLXqLBP8h9rqzKaEfIJmrrU5FHnu2nmwBe22YameMIfhEHcrq0ALDRI
ZRo145Z5fBykTBZYQ2DQD3h0ik5hDdP56GXfuR6ceBFZVdoNcEOwiwYGHsZNYgVikihR/7yJJBYh
twqprNpUMbwMt3DNk2GlOXiqcJXN0sMXMfZg3wZ5AOkq/dEnyTsQYFqvhb/QWItIUp6+pGoVGUlH
bslPuGVIidjB9QQu/n+EUc7/0RrhIg+zzcnRo2DcB5gnw0wKa+RoWh5uZDySMwpX3JSvJkZGQ6K0
UeiLXWeoN/KVDVF1u6o2nRzTU1tDFRLc/4wowaWjRJO8HgoMLvoZwLk/7HLE4JU9yvp5oe8+VZiE
zhPXwLC/aKyzLs8CBCtquGlqpbZHhqvX75yUaIe1F1tlULQhoZchwPyLawhBd1/yI0/WO9LkEkra
WHmiizWa4jH+GByKd6cV40UID4ypqD8BuE6FKVYfKGV7fAakhgXUTe9JLcCX12n31+oSE5Cv9/Hc
WMbx1isbng9VTgSCCF0+meodhjIPZZdnBMa9Uo1szjOGvvC8zIpouh/ofGJTGh2s/sLAHhVXiWqT
Z4+InUTAyya6XZiwlRv1AK+xGTW9sbYPmEjzZ4RzuJH2Wf4DPj3erqTyYE0IRGZDrYt3KdlGnMsE
c4+Dy/iewbSQmlt1llr96xl7jgs+bvdoB3SlovPS64v4lKXPju+2E6oAPpE/26QoJTWNEwVpfCqT
LzFsmnecWTli/O17BTawBlgY3zazTIEAF7Z/XfDcCn4q9REdesYjwlzZGB3U6sw+o0iv6+o4Dn99
27WaGQB/7eLB+x5mkU/vvCeF82oMcJMtvj2CURDTHOY3V2pJYPxJ5wB87LzjKmW8vxZWch33doGw
Wx/wa7HfwINVO8PaJYerfxSmbiyXVZcOOIz7A95frboCHH+7DWmCAp8KwJuvochg8w5DldNx4oSr
E9KhaAga0st/eYEnbscLbhtoHxD6f5QXi2br7+DyY6B+bIMvYhhrozYizljn6a2TzjlQecmFrgTu
odgnQb1hQoJl8m8RwRdKkJuNw8T7Ka+Cw1Hew1oAsuyeuqtVzA18C3HaIFVwnyfxQfiiHteNTU/X
Wic+vEtoOaOFTN6VeVjzFk/ipUBBkVK6jphlnaTo3ZpoTWK6yXfHbgzlJ39+L7TP8JqBybbGAp9A
H+QsQMSu8shfHq/emvkn7QOzFhQ6WQur8LLl/Tot7xJiegcPSQkdlIU4ZxQyrFk8up/SDGxXcbvA
4/KiVdekhCE4Kiz5Y0w16J2OKfm2HhCjX1bHDeo4DR+f3I64dtiXbque9LlTiSXFB+Dn8UCWyH/s
AyTfootB4fMiMb9sTdk/xCc7+zB2RsVDeHZeeXcEG9MAXxKNxr7NFh3N2u3w8pjLVnuapVZP3Lrp
5v3qZAm/dtH3HkvKZNyYyTS2LgOHipD7i0qSZO2GiNThzx9g9ZvcdHaGGffkPUF6RpS2R4SQ8ccA
edWBY/wHkB9bnKbvyTlALXE+3XeOa2eMS8j9PhCw4uVePhSuf3Rwy2iJuyYrUZWf5BfdvWDN/ovF
tOMTrLkVNTWipbfgBeYCCj1M/A7GqJmZ/53trj/qZibY6N+dGg+mraH2uS1NAa5eb0W7vQVjoQ++
Mxx+frUKh3bffp6X9GRnRxwpq3KBJaltV/34PWDsqMZ3wksXA2Z+a4NQMxITklXTQKW5uFPirQPy
cRPtEyVAD/eOQSRsg8/5NZ1w972Y3czHTA/SrLb3TG4QK/KFUlsiouuPYf5G0suEo7vd3TeGpPaI
n6/EsQDm9eBxx0QLuNdmDLDQe/Xh++bdu8wNY8X8XW4qM1KfHZxW6O7qGemKQMFS/9Nha/zkFizN
RJlf6dAFjusH+vfnc1g5sE+GvAMTV8ElQvXNxMKVH8RdCya7vYgtCnSKnRLo+uTMyX3m6iySnGtH
cj6/wrF3b64/3+rVpX6cp8jGi9V+96iI4yq8wmggh6L6T576qrA0Ri40udFWMZUpQhlIEAEuHQ0j
kQi7/IM14Bpaiz8/zFy2IiluwOZJmKERSANp4JFiorPf3AJXY6TPwOhBwvAJfbQQGzIaAvNNh/f+
qWmTfGjCKbltQdT9w+lwGnAXHl7e6NbZsOJfjnrpMR/XN+UoqES4anvsTKTq1Ca4v1CkJRAIaooj
iejqpCcMOXA+vqsUR8Clw3c6euZeT/sxPcNTwjWX80vylpGhh3Y2xaOXu+931ucyxHQki58vOAVK
3rdcf7p9i3h1HyD0EBMKy226vwJcBwFoZ/8b+LPE3dpjaP6tUbByAOTHIyC9/AXHGe7yMTg37dBQ
GDC0ZZ8TE5nV6X5CSnDGRdXHOHNsB+JHmGELmdhW9cknyXTT+WkuJVoiuLY82It0PcthYa46aN0E
1lYa1XQQvpauEsTPOLP4H6/oIdIIJKzmSmABelXfRLH7toT+XnLI3jDBbCp0ynNfNblWRb0PeDP0
BH1DipDxKeZo1mQ9tkCIHiL3vF4ZO8qyWalbklPZUdrAVrVrILYgBFm3fyb+ZmIgtuCx39ImDgJQ
Ro2wmKBQlLJHmaPke1jWqY6AncsFW6y57Ss4f3md8H2V4GY54xnzBpvQ5zNIgYo4Z4aTNDVaGhi3
x2tigPpnX4gvnjzTNrZnajcJSm89xzjNOrljPY+PadjqSOtsUz8nQX2H1PcAVj6EQbaH48M9NPIi
pvL+NmrsgFKhszdlyQ25Dn5KB+Mbpy7YTfAWF7wYKof8Qq7jiGlTkAT9Bqk3CQTd3Ys2E2bsI3rk
8Fe65vq5dZJmmoemEbxxWDvWjtCrmfjA7918/HcUs291Gm8mYHLDduNeAeBdCTWYGIVSdD5zm128
BvUtwk4+Am+e49xPSb8EOmmjTg8Y/C0T54o1bV633vAZ4PXau++oH2iOr5ZKIoxdbfFLsEo2qTTw
OHlMO8U7f4T4/2xbUNeE2T3B+TQeDUaODed8vLG1U67+vV0AfF5SGDmmuQA1Bv+P/8LYnugFEPt7
F1TzwmwjElZZAAxKUcCHGA05GhkCaZYoFBO4gCOhA/KKVFbR3XgjUgV7sfzByslk99hX/YIZEuu9
y+rnww3bHKtFyJs+dtI9YyMJ5CAUiXRfI0mmBU4JU66aXsi6j9uwV8U945PvBZAuvnvTEnwwHknR
htKBI4lGMBHUlCWXuWs07Vn9h31O1Yk4k8LBHYemQ5T02o0SpWdFQ1Z+4MPnuzluOKuwZ/7l20PN
RwRZDZuweG8/0yczfT7CdLvJOHkOEojy6e+vCP5oK/4Qm69tdVUnJ5230/AdD2amfJdk8ztr1/Tb
Hwiuko6bAoK1ncr4EDxod7028UbJ/WhWq2P+kwiElC1C9FgMJ9qyCBQz27fChCAEUMpr5uAP6gKk
CJ+YYJcyjlyJ7Mhowmgqeee8dQWRpayXFX+/gYo+t6i29ntFfBDg1f4O8GQBpaQhlGxeCjko8Wsq
1fTbKPHJR8KgTAcL5wr5QkUcRvHJ+BDpsI4zfJkRp4U6zzrS5pZ4YdaRnh1K2yppt9ddxPpH7OIF
oJiWGcjust/KJu97V7Kc/mlC+5Pr0B9qn2ij+0KOZyalQXg10sLfDptOwlmwWtLQFrCcCA5b0z4t
Ps7ymV+vcIe3Da6nIMOvSIzzqyeqQ7BFvby36DEE+BuOfji4UlmNmAPgqDvzc3PwwV1xQPm/+iYj
GiEcSPgOZdJHC5LNQHnfovFgzIY0xqJGY+mU+o2JJEHSItAhBNgPfJrJwONGHqdEnM4Pu3xjIuR9
AdTyc7RFpj8qeWF7ZDZj4lQuIQXt45ZyPvZ/8y4+/8lzIeftbxCfyhUTnvzRnNQIeAKX2YdiTYAS
tkdY8yFLXDRZlnnzxOqMcZst3sYoTauxb3icdu1jtonypWAFOA/WNoAZq5cFv7SG0xuXdPdzpdbd
b/lLXOBhfC9RqmTzWySxZ3r+dgep9mUeD9hjOr0gD2i+SRyk1qO6IbfLm7HM+NVDNrhBBwvA6t6A
Ywh+LXgQj162/fUGj5FviTV4QqINwaESCE4jVNZL0jIQ2Nogu+Ntzm+f5MLmEsUdZmYYm3gjNBkO
csbhwTUT17TfWxxsF+7TUKwnRWgs4/k3UFEwhyZEYPzNzXaowSmMFO48m61y0ShLDsGhxPaehH1r
nACk/am9GyH2yfvG09yKw8wcb/DCdnIlUayx4XNTBV0UH7MzFsJIKBpfrLU9ixq08ubERK71aIJQ
nxScdPNzXpSjkmAv3U2Qhx8Lrwantiptnzzl6qV+tP/ibdjDBfIpvEU4foVDcSRrHCnzAMnQKJmn
iQwkzCdgpyXUUY9996OajtuaHYnxrakcU06eFfdPHfqTWP9gR+0bYnsbSFWM4kQPyDNDArgq8dRp
1o9wXwKCCMv1A/ZZY7qkWbNktWqenKteia78Bl+V3BGYGdC7oWZeBEDnVfek07jamCpTdacKQ8mo
sZJ2dcGRAUradXkxYR8urLZxGjHkTuw85j9tqj4STTWlaKhv9Z7BFWEIEbXiusHmqpPlIkT89MJO
vbcrW+TBCG4LE4DaCbF73/o+vUvFLFZKiutx/zGmAyeV1bN/oriP5HxodT5dZOXXVLb4gAYvD+xo
82jVWiuGrn0Q6PvuQMAato2cyEV0t55JdniidxhndJdWVJfWRIeJ3yEspOsbPYTSU55zQgRleXA4
i5f5hMEN+LmUexQWLpPVxaTIllv34Qnli2GbnrLcmAwfXwtrao4wnoy5HZ8QfDxXQOkCDPR8jm4I
ymaPq0JsakqjP8syRLVrxKFzp/51qPzuGOgyHDi5ni1hw/elSWX0XZti8d9iHxPFN8q6I13rGcmQ
6NK5R/Rwv136mXbDd+MhgjfbQ+KbwVqEClDqkHhS00szNXBYoU3Gmka1JcnhuJ2AanvnoRFTtdx8
4Onx6F61IXpyqFV8VLCVKKsT0Xjn9rjqlTzB0exZznZXD0WYE03T2QSeCj5+csCG7NriER3SCUXg
DwsRc+k36YanlTL3Gt8OsO711t1CdoVoeKdtO3NFjXdRFEEOZadcsi2vo27nVZL9hsMkznBuT6aT
/XU3bfCFewjuqzlAu+QecX5H8KgnC0WWvYWvJaoTxvZLXql7j4xSj5SVIPNOr/vmpugzb779r26i
9AAsSj56vjlvq46kctM178nxCqpexVBLgCeZv0b06Da7AfVDXFv1MwlfhCfOSVYvGuI+yWBNTUwO
SFLpU2E9I2BvlQVlkpUSLEsGVSO2zboNXrMDKtWuG7Ekwog4iE6rZP4Sp0ffxt1tEEPQwudGxAb7
IY0P7OZmLIKSLWsxOv86QjyjGaxoP0y8kTI8+JbLPY9W3xLDQWF8tpPY7+7fs/AAyPlo/JCHDoFP
vFd1+A1yz6urvQ+MMCJWl+pdxVHqm9uSZui5w3KRIFvcHsi4Rp+kQdeptbskoOqAcvvQsTemlpWh
JVqc+H89xSWZlRh1KZt7VtMmADYbalEWYPBmzVBUpkRrHs2tOg98OfYT0X/o2YpN9FiHWnTxWaGQ
k7qaCj2Z25XSHxgxZ71fZmR+UQi8E1tAbEmI9UwtXZZH/IGS9OOBTxMgpd6oaQ7vD0qOx5Uk0ftG
Fip2KLOVi6rPWNDXaffcn8PvrtMmYWUnuFa3n2SssdYv/QFmul4RssMzlPUCc0kytFTbf1RXfjpb
8X4kdWntYmPEU1muvI4681DyKjpr8zvGq57504Ww0cNIoknoOhrcj5GQ02m7ZwkiClBsWBWmwey7
yJh44TV2yucmmTXt4UKEZ8qdl7ei+KRrv2m8//cdaGyagC4LMufZ2frNGkdPIrvpB9vYE3h2Defh
l8P2gY3eiqOL7uUfHabskmK/iHhxF8179/GQL1hpt8DnpshDa2vFQFb5rXJvxg/PJ9h7bNy42L5K
5e3RO1D3cDYVnZlIhdN/THBe/MYFPBZfGo5diXovsEpfrUrG2m5sp4MIK7pGzsJeH2dB2X4oC3Zn
V8k8R8fJG52ppcdRimG6DhtznFrTnO5FXQjHHXMYO1H/fBtMlr1jeyGGYPUZfJ74WoI2fHjYaBjo
Hw2ZWXXrhIrWrqiltD8JgfgXn7Racc7sYzV9sfpGNiLrWqBk/aJNR5hnpHcgB5k3btDaqhgkTC4H
QBjCXGa5O5TzKsg+h28uGNgVX2vAf+YewhhffjnsjJFmsWcl/OOla8SfEG9Al8RG4/Q3RYqywL5L
2Xy3cgkfPTIHRocwmxSVWyVcDcA0z9Ni6FgvVMrrBTzB1Puab02sw3irLZY+noNW2qsQ8foCAlpg
7gk+xvAuzwUUNaqLEIKfdr9nxRzMp1ZKXOXpJ1QD6PDui7hv/2HmXIJRYX1sVsoF6UROTyMAu7cb
7lBaVXkekuciSPNojEOQagF2yOBnklhTHmDsJfSxDRs7ktX1EAHgEHx/Q4jcl/74FfWRU5DZ0s+c
iVp2O1oph+MrTAp8WxfBOBZXrlbKEGER7tJe95pE89IHGG0g1NNmGzuqNd6JtdXR2emyQP+PQnjQ
tz01h4XEjfajWrYqH6zqR1PVkTGpvV/WROX2n72YhUkCz+6msAad3LtBqQmJMxZMypU6r5hbnmmz
kIgHdr0QF5TbuKn+6ISWXJaPKIao+A0IIDKjuzjv5TMslNCIiarFyWggcqO5XAndIyhl4BTxyESN
BLCxs+zXwH0/FcbxiYLHXXSLC/nYAJylYSdKNl3HrjPlMNO+FPFKc1Q3z7cAmkI2KvbdSMMs26id
HLp3mL9QTB+F0DFnVbtSyxUe/Imlu+j2f2gfgS6UhGYnp9FxmIFAusRmETXLr5z7swUkNnKbcZl9
bPSbZb+nkTlPfzusb+dxz3UCsBaprajHtoqa2Df/aom5iF8K50m9pTn4OolSiwf/TkYThJ3vJgsA
AGDDUUDBm2mCJ1EzP0U8Mq3Fkrl+fn15KfI6zjFrKzZZWGgayFrswT9vSFe04xkp47V8x5kZ/soQ
dSmRRW3o5myfpnIHeLuHDs/x5WQQ58sUggF0N3kEiGRK/qVfW0x6mjxJavrlVNTU5FJnQlAs2zLz
FcEUWy7OUzngYbaYKpTCH6uzwaBB+MWfCAQnUbkLukRo36cz22p8NDjeKxUa1TuvFENTl9yBZBjS
ic0irrP3Cjfwg2wgpH0evaJjBnC8n457pZrRjmUOGJXHu8J2m9DMyX+K+K38Ps8gX2MvSw46d7S1
UW3Ducu3ZHtGAaubky4Cgqjd6DzN67lHs7stCxpo+nn62QOBgr2pURlRc/MoBp/11/H2nrB0SclM
+zxeVb9XiLCPspc/suTxWE0VwUMhluo0lDpcPcHYvnD+M//b4CDZvueL4fZ1dGLositTcFhUdaD/
4+uaNjYX8jHbmcpQIJE/vTlBgNpH4KVn7/BvlZhIzBXmCrw159mQs5bniVm1DiDfR+1tauSBmD7o
GcvxU6iHcFl/sCtXDbZeLJ5ReqmO4KdExfLekzJBb3zOLVBHxrNRV9xM6fWPr0XFZ4sWscQ1Qwjl
YIw04DQUwMegWH6p+48yxebLMjLKPC7XF2ylhEYsdgy1aLym+bKw+bA+Taxw2rL3G4N8c2z/B9IH
AnX+pxeP2ejRn6e0TJwq7V34aCepimzSe9PtfvZX7+SHI+oi/OOwMSj5kgtPJnGvknrEpxCYivO2
Dw6SvDq/ONsu1O2df1Dex2cikdI+33Y7ZjVk8QmIps7wvP69fTQkGnywksjUBDsdeQy05deHOVF3
tIz3sWKlUSWpYN3c2OnAzy/MtZbRTN5Dy8OnGA5ZmOM8CdAFBrwJ+uDlYr/FwbwxDzcRlnT7KTw6
xs19Sea+GzfOQslzaiTHUgUqg8QKg0+qMBMbBFTmBkQ5ujXN8RLQuYBDiy2jyIy1AxwbnDHgGLcu
wKFxjtinGv3dYok1DylyFVBHffgno6OA0/eXT2UzojjsCsBBzmtmyZPAakwRSLHYzO57cMevCx/X
yTgJ7Pnd7T/kRkUCA0sR83FWV/DbeDtiK3x96P1O+bkgbAcSxsNnCSETVB1xzzXiUMwDQ7F9pCwf
i5rZEEB6SlUU98ve4L0Zhvh+LKVtrs+YkGuO7kvWunVtsOGElx4kUt71NF8EcIYZ55AEPxUC3hf6
Z7YiTTAyU57jZeE7fuWZ3b26TP8rg/Rhq1heaRW8U27q7jMmNFv5gATP6Lk6DIaFc9GYjZcNsU7F
J2ob2fRCe+sOJBOS4RKvuhcmlxBvDjEfgabODDnKpjS5GqGT8aj6AJHcQ9DnO1Qf3RYfvHL2cGkn
J8M2uhwd7U4jFEewt79bVWFq7KlkyyIa77qDLSggAj1sO2ul8qaXHeKCO/cD5D/RqDQDNSCK5MoZ
+PHB/wcIar1NZcsV1nzOLvWcmeZY493zvYP5VUl9lxzG+NQqp5JCo7q1VHWHAi2NY716T7h1d0eJ
9o1rttaG161RDMGQFoQbU2ptiGsa9CggiPSSLMGuxum54O3OfPZbHaEpASVctUnyXkhpTezTc9Ad
HMzbxIAA9gCMkTKT/mg8LM2EWJyzaiL/r8QF6QA8ZjXWa4D1hlSqiIAJGTVAEQzok0eh8tyM6O+3
F3sSMBNWUGHcK07M2ywCkqY1f8fMfqFA8tDBbQsT+V8bSI0LWeyYguT/LetI7T8MZh0vilxU1G3A
N01HNaVJDQn49e6Ca0ILH2TVN7iCaSuL/Hb+tsn0Hh4hvSZpK3H0m74tbRooqOLAmATp7oasHtZS
F5VwOX9jz3VhNuRPYAcRMh3LcCjHFc94DdUJuY1eAGNpBgTu6HvlAAiSBsmViAi2y3EIzzGY1hxc
yNV4c7gh8HrcYHOioM2J+RQRw2Kindv/fuQGcgDKf6sjclUirB9LKzMfTj5Mv/KhLNPgdGVUuFaH
qjzhrwltC9DWAix+TYt0qbVVezNjLyJM6tBi1ujA2EcXze5QFhNaz+ztdfUwVrg1lz0+E0F64lye
i6B/Wxc/I4SST8wlsPGOJI2Fp6QGVFFV3uAotg2jKvkPpknXXc++wzVoGl5Via3w7wLvzkBPPsnp
nfFSSMgB5fxhe1H13rdycbCIKVldKC8mLulzEy2VKI+9gF7dDn3pdh/DdPWqXPP+bGryDIvhDbWi
gUofruGtnivJVfuWueVIOIxpptoQB480WfTiFz5ef8nu98U/aVkxoFs5OtU1M85dPt6oD2DAFG1y
HgcRcLc/QfOoC7ksJE44kwaTHGnQeWWI6HQkh7CLPeUzK4qJ4LbABm3KtPyIY8aAFmOOKFqIBm0S
qnmKDqarDuczUcJOO9p9TQxfoU7M0XTYuZohvGN2a/vEInN2rAxQIMtJBsUsxBnSqHtc8PsGQC7u
3lVE6f4qGdLTDoU8gm2MrQAJCv4kgZOSL+l6R3Bjb2JGnSl8mWbkfg/iGYe6gKAHd6QunHktVy7n
AtxAva+vtqcOoVLOa6AN0y9y9jA6yVXJ+pAGSdkyvXa5xECOf6dwGE1xuDrKSy6hryxN+hLqJwT1
rXiGUTaSqFjffwxuDpli13NaeiD4z4+ZcDJQEWomGJwV6q/RtN/2abg/FSKpbPpBem7ZO0sJ4Orr
LGEPywuyNAwzhhMdLjNNj1x13BSzVf1XmF4TgxBVeK/6KwtW+Le8d4Urb/0+E9AuMnV/RQ6N9vRg
GuqYec6H+U//nX5GkQ6nckzJUEOVnkB+uAeM4s8zYWlDk9zziC0j39C0VcMlGNxpBaP6mtu3NFqq
TANqdta6UjXfs/NZB08qd3l+SbdjYqS0hbE/tf+m5LHGZGbtGJtqxpGOpSnO7kZZVDV+7+YHb+9P
e7H5ZRlmoul9aT+4I86s5MBxJA7T1is+95IjZB5zB6TRKioxwq1O0e/NEfXQBJvtj7Ogm0MRWzCr
LCG/4P0c4jqHrWBYLmE+fQsNvMDqhygMDVkb+hoCv3qPX7/SPwGx8oalKF8Doau0d/aetYxFgmsd
GyXv0692stAmOreQcMQQu/sCcwR56a81lUWzDkNXFGtbHPNA+zxt6wdsyRW/f1ovuz1boEPkL7ou
+JLw9jw+FvigYeXPMG5B16Xx8d+zSCtH1i8hs7Ak/Smhl3Kb+uHV77wjpuiyTipN6//HLRLW2Rax
1hVEyRBEQBtH6iP+ymMneELdjXv+lwEgDpYbGTwzs2YJw3sOnilRb8bNXTU5s4DhV86a6SlQKPXT
jLSXZ/xBC8fVLfoYLwR2xVfc+1bli/nyjV/PelAMjcJYjZSWmxdBe5fOOHvLaN6NnAnL4CASEgCW
cC1dAD3k0YKadvdThNayNDHYNxMSjm97Y+8O2mEYULnuTTsuniPJFnje36vqxEW6+ZtmLdCSsSeA
ZQyBQc67RMR2f5+/eelY2sKIIQZMGwTuw7DRtEF26HTaliHR3EEobnyqX5X3kxb9SDCT1p9bEfdX
qm0UexP2xOOlwptThkfylopzfFOVYdn5hc7IfL08jiETD3QnkYtc6nuQICkpnrDub2+s794BTPtA
IAbA3z6fu4LeDKZB8a0qhPia0Inh9q1jaxV15/BD9mecSruezKCZRGnTwlYcvVyxbFPbT9tIERHp
1HygBpKNvzbZfSPz0AQbhZpLh3kvD0OWXxTRX0obDnmc3/+dzBogoQ6YrICNQuq9C6oQSNF3KEDe
jLC+7xANc5dEwYOKZWDTT3f4YKUcdYn3X6ux1TPwqAsoqG2L5itWB3TPS+2mVuhBfS9w8PgEHkEz
MoWSTC3BsxwP8X4R8ayH562M88axaZZ/yMl1KqPIc+wnUW3NvtYB9LRrk8jUfu+tU5sL9MKbTGcb
Ij0PTN2aUOq/BNYxbUtWuqQJHv0e7ns0gy5Lln17GdpEWWKQYZk3p1M4bUshL2OwpGW6j0r+BB5u
HQf1Syz8S8Wmx3m3aEd0UZOkleqrIzMSbqzjIRejJWixz6Q/YiEm1Q8/bVbJjA802+xFlmyeff6N
XGTD/I3RlQEllFBfsudiReSXYzIGUE6K83Ai8C+KxF5ywlwrg5usQyCnZ5Pz6UtHx1V4/M+gZMh/
tnuUHdipbXdYz6neWxKEX6vIr3FzrAD6Q2AuOb0BLtS9bogkKTAfkFKhGX2flKVErLiJeXBZvDW/
ixld9OYjZhzLcWrjU7d75x5OyFgFhqoBQVFVI2TDXeNAR6InDOq8+61Qja4RMQTn3gZjyonkY9UM
CLn79bCDGcmDcnR5Vd/DEAkaPtOL8aGTgr0ys2rHYCySlUbPuuBkvz3I3f06CNYsZfVVCYcXpLIB
t4zqCK4W222/otL9a/lLKaFNVh8XL661pLSnHM/0iK58MpRFexbrU+xTmA6twIq4sS6q/lWqa+Co
athk1upujYJDAYj8nrp+4A8bk0p+oe+257svmZYxSPt4jNQMSIPImu65FLZsd5nUEgSrfLbhB9iO
bQ21AvvXP6pUdpwWTpgfclrvyepv//Fd+LJ1WfwowLWEkKPQQEaiZnLhA748pY7hWyH1Rxc0p354
hJw119mNqoZpYB3MZyr0fx73d/wZDFs78ckBIwLGpcyUj2bAyS5+5mZVcE3Mt+4AcO8rmBCgy7R/
ztVkxuV+5vzrbLktebuQZZHocmpRXeW38aLgT7O+PtZO7bVKouZkaq+UOdmKwc7LxWtfrFw7SZU4
nIHtpMwssAXMsEbDij9Qap4HTgCJwinqfi0KqPw+Mm9nfrHVH+GG2LKDt49gtS2QUagxmXOlL7k8
LTtbP9PCkUA0dD+3p481tAXizX6dkzwIiwq9ZXkDu48XC03JzRoJWpU35ZZmkmv2D4Io2hAra6uV
rrZ6cmaRCcapOw6BXaRXIcdgQuuXp0g48JvLSfwVBUslkA9eNZdcn88S5oqbiX3pWQHSMI4FG4pk
TsERhGyhdvjwti2mmrwwPfuPRrtUqGZdly0dNTqL5Vo1A5b5RdbLokTGK0HNYuBE/RrRkHJKogRR
2q3S+oNiWyJxHbYgJD2d5t3xiwao0ioZdLeRlt2bQvlfmPdsY839Tap6rPaWzI+M0VVbzYi+0cd0
+jzdEpcvjGxvQd41UdW8t9PlZc4gHF+Z0wAh6ajGNhbuBkwIkgxwyBOF2gCv8+BSF2otuxHmsWmt
Y/6p7N8DwEpSnJFx363UCRI/REnjRgBc0wi2Fp4VpNikOFjp84Fk7K05K8tm+XNd59AIkbCt4Oor
1PE0ft6zii/Xer99ccYOY6hfjVOVXeHFLnIi2kbtoBnbLeZ6G0rhjyp/XQdGSUkzE3smoXGADT80
ilYdsQU+/rPzfKf6DhowB+hOg4nUa35FkoAaOJhSIvqCeWGoVEPlNkAO4ec97sJE0oYHVm6rbk2H
yGdWGzEo0FOWge0Rfc1XOI5y1XewAcDUs92ZuP5TyJsqQlJVfwll00mvt64kY6M+6sbl+QdS9hP/
sDl37p8sSIvRC9tioV5Ap2kw9xqf3zjbGTWsWXc3luHcA6y1tSqnd4pCURZGhUuXFm3Fv4BheaAF
Y/FZQizpoa6txCluJRVMfiWcOMHRJo60hPn1nChzEH4a3xwypVUhAiUsskBUFC5M+MIA7Phw90V4
YI8GU85AWlc9xzjRkIoSwLmDeJ2lnNIBYJ16Suz/ItKoUxaDVg0kXPFMt4RYhzTwTAZ+zIimO8h5
1UaDHosHdC34XjSR7H0e8nVt6WVpDc5jXM/etZPNDgxMX/1OabLh35JOgBjAFjt66ZqDGi+xDHMm
Bf1+RljAsVJw/2QUYnx0FVimHnp0DJhCtoDnvv+MTCp0vdaSBMYW1L3p7YJ0KZNnIt+835F8z1Uk
Ske1Cq3gRCKofGQ9rN3rE/w0ZTXPcs9sIP+eGn0VLffLkKEP2bwshQXoRMJNHaXkwL6x4LUEtZXD
Y5przCYzDfzW7SdMkvqxreISys4rc0SRktwk+AEvZxWdi3zm7EN7vJjc8S8sSiOnGvVw9hxIp7mU
G8uHxQclnV1klGygA0lBhxlaZRrL47TiAKGB0C5omNdlNF/5XKdw9e8F96YEzIWV9FnLVVYBwhtH
I50y4uOvD+9TWWWb2m+l+uJlRdcYOCwH1DHBTDUyWNbHsFw+lZul8wD2UUQGUY86xN5Xw/mI9g7/
qfLvht10PWuZpzlcq4KDOb6TK82UUWWLw4OL0gADdw4PE3fhXnifPuCc7ca5oOe55tnnBL8NI7t5
iHOXLaIEHrI+3eN7HkitAhqhV/8dmT3h1cda3I/j4e3nBqVGpQKhouaNWhdfRqB4rHBiFzw3HAqx
UyMdsi0qrwo0c0XrNbH6V6veQ9ttLx3ezM+CzYmRGeqOgLLz6E6X5HNAMOGZZP10ZRm6ocDSY4qX
aiaHTSuWwG9tZQKErm65/xwaK7TPmYvgKqYUdIRI5p2D6NlrVz7QhJJBXwggAkJSrXC2TjySMaoc
hUG9T1iCPt1cHkxN9MqfOcRpZ5YDpr0fX/gPg9oHB4QcOKZ8UWIk1Pr+PVhDiGI1kVutJXuvhqVk
qTg27HWNjbRgqKXgb4XAV+i3gFe0a9TkSzimVU2X+XHq68YtNuJq3obAMuRdyeOtuDFptW7PMBuC
sCb5mL0QWj+saSPkttV8sOYQ3k4Ldd/nuYD8mubMqcRwH2F7kyTh6/+KPp9tBlD8ipGDAhUdOQF2
d59hTkr92M6zu7/Tc9KsQRRwQgkSi6mBRaVldMquVfFq37VUkBK2cfAMh+fBTtzGuv+dwxG6GOaa
GT84NbcWOSy5Em9IEsg61RgNdvZERx45FxDI/H9xYjVNYr4LWw5CK5hNxEvwkPNt+78yGyWf6FPG
PWGFlxeJcI7ogutHIzCZbjZQ8624gvBqKTgawzf/PtpJlovvHZFKS/Z++pSdQRKDV8EPLOeAk78K
c0PwpOQZQKcq+R6z6j6dpt5NKLcu9uruehJHN7t6MJ+aOf2ZeizqappEy9ZT4sMTwDWHc8JHvV+w
UPuOsBMQhZ+Cvhbui9fpce6loQgCgTqRVxk63QfBGCmZ6L2doG56ypUYu0kqw6np4oehRsAy4qEW
ozdUev0YUUtbWeutijM1E1dZKznBN/pNPj1uLBjYI5J2H2T39p625tCDTQm3y1Rp8uPOIDHI944S
oF1CAoOfe1HyhdHd8ShbIbmcT8f6g/vB2O5zjhgiMxpcmo6cp7V+20ze0R8ier9HurAs1JhYozVc
OBfoa8Lkf8VAX7ReV3fzz2tJAxTpRsUQZGJ23ngj2qKFEnZ6JvIJi1dhgOjDypRAiTLUNu2wov5G
MflneakIQfpxYIAbCRurmgcD5fJlrVzi/bcUMH/qiFheKQwdEQ7HLzAwNmbs26I6dqeMnBaZ8aqY
uZ8TLHX/lc0PnRC37Hu8gIj/rVFpQyf0YGStpqAssVuGRoT91bn4sn01jJuNEP3J4ojdKXdDYOfT
RE+OUqsxlTU1eQl4989i3KMHkvog2EaigsgAXyPAW7BUM5EavHlEZuH5+DUv4aIBwhIkUAG9ZyH9
YM34a4O5AGq2/m/bumvMEGBn9yvclOZN2WFWfbLP3JLr8zjMmnieO4sCzXI93HZZYSywclE9u6fp
THTs8a6bGyLGzcCxnuraDZe3nLElS+hnhoV/BQwkVAZgbn2itMDDA/5eIlMSoSW1kK5zCkjFayjy
cq3z89obQDO0vWdwToHM435ZS8dZRNBQSujnpyRGGwCUn2vZDvXt4oAthGvDjqc9dzvzxdGMQZLn
a2CJv0259xU2++hzrNIct+HxeqdYgGDWAvw40ScL6hHAw2UcSypvpTCxeAmlxDcri7vDzRQAd9z8
ugOjxosoty95YvFqWY8EKq1GWG+uu6IH0a3GRG9hp2B4Vik2ZiJtMT1qBUkGE7ol+FCUbPZNmL7T
K4Lb3I1I6uO8RDH7sELmWbfdBi87fhrYGnickTmgcWTpd/sji+lZUibc8q4mHKZcRJq/UR4kFJUB
6IzsAtRS4g4ZLocxiLsUBHloJ8zFs2Lp9OfqpueBvs3XtswBQIs0elcIotvzYB/VFiFYytonnsBC
ra1xzO7OrOdc8pNm12Yd+j0CZKqgMn3lXTBBhu/yH4cHOUswfTG26pmnmyAYqrbj9yj+v2jUNUGX
/BkUXyVqAZaFdfwhbptQvz7WOv+qgOU2zova7FMF9eBrhz+/2LDgZceFW2NP+gcmVuQtODatEDTf
1rl68RiFnlSwDpPPQsSM1+XMArshrMApDZVjuHX32cdOUBoNykKkG5Nwq3gXAfxrKU9vb89cEqF/
5neonqmKZvADO/xc8FJs0LzufHlCICneDzvieod9acqWKgT5wa7g+Gc2/U8w/68qpL77rqc2B+S2
Q2hTRwE/yNl+Dra0I6AzQVzAwoH/GT1+wmzjxbAADcF8qNUrgyuB5ZwM3VO5OWntRcX+C+JHfh44
WR25KZWSsI0QLcg4M06l6yBp6k/qZZXT8OqqO3RmBJPzaHbyRQyvK0vf9zxgYC+FRDLE1Yh8ZciK
PjtEzqtkt7CW8HwMaE+Bq7a+oAVBKOwVZ3toq8CtpSRUhfvuvwLCkBEWPKCO+rA8yRl8GRmTnoqL
HyrgDaYX/Ob96/kJM4GlrbpGQb0HuqVN78/fFQvjGqECB2I1kroqUN3aFljUxSsGu7TWst2ozrs4
VVVYkTLfmM8FZZ9j7iNt6JKKHarWanUodKamoWOWkDUhZqvlfVvCrHQG6BDpnyCHKVKq9hPuG8a3
QV2/bvucvCEEYhc+koDayCSo2Lpwbc3RGJQq37vQthJOpLN7g/59dWmS8YeeQ3kIGXZ1l3a6nyo+
+QpFmXutS0TNWCe+xYa+pZI+JXLbhXPp/2NPpseE6o5DVqtTuerk+chZfn7JvGuxTXGU4avg1HS8
1f6k4gApG1TjxTyLYgbUKQvHAm8DtChYf0CROTRVNtx3PrcpPuLe6p+tpoEBmO3g2SoWHPS782Ct
l+nulSkspZZWDdz0VSL8/tGU9YovmGwwx1rVbGN6fHql4l4pH95/7uhC5IyWwTxxG5Gp3P3tFJpI
Zhoqt6k4X4t6twddgkyzPtrnFLxhqDa/DMu4n1mYywwBnFZ3bNtvw8tvvc768ApSU8eQcTo6KlJw
mwRAjDkZvGEBBaYk5d7f6ebTbrOxHpoPRlG2aO4zU6HYPp2ttX13AjZKlQca55k7cMEPOeBbj3OR
XRLBFS1lgrZPvKYvYCCY6uDaZXpvXDC3VC6npzgXFvIfzBtai2NULlah29iuSyGAlbt+d9ZzJOzb
/rMbwW213qEFxEf+pafvIS2zYbFU98BbquSmK7R/fl2jMZBJ4YqrOC/FUZcxy5GvbIuoA6Ie5WTy
DqwSpg5JmkHw/lDK+AbWS2DDTzr9MtMgISDAH+ssk7MwHoirJCzdpg+6RJKPpGV3SoA172YwGakE
pcG+dMc3VIra/jmi/grwZ0LFAzaJsy0npkdunyQ/m4EDoFB5gkBtGQIPy0ZrH8ze108xQnPqTzBw
uvWmFYnU+cLTiNoIUVCGwlg9saHFD4q1xpTu/OY2WoraFEfmJqADNG4if5vbSjeXMl/OoB5MkIs4
QMLdOfZ4GN4E0BgdMbNLU45sraxZjGeTh+RBLNwiIkShjItmTT+QLBWPg+7tNzmm4rXZKUjNUXQk
qqQVTsE4Y+skaMDsjzyBQCrB97YR2WRPgp1TBM/+h8CC88gZ0ZwU9P2BSee4SFk6CRI0HmJbiY5X
3ToLvgAI3fNi/jKMkI4C+Hwdogqr3+RiK7EUXRm0bzzMrIZr9BFHS3skT/Q2aDb0VuXV7QVn5VS8
Q9kGWF2bi2W3GkrD/MN0mKoU07GA9U/tQoPzRLjTQgToTf/8N1owvBG8wQ89pD/Vxy5k3RJKNwYa
RlGHBF5on5Pwt/amXVpt1qG2dLaxeyd6fKWrzkPBcA4YmZyGhXA+NP2zHVRedb8Jya5kaKFMeUXM
Iq4OtCd3jdC0wI6zwLr/deikMwimlY1PGqyFp+glRnHiYF1ZwMpuAM4Tzj/7RDd1A6N/At64TIOU
Ue4ipAv8HevbOpo4GKGUxNjks8ovbSRfiHX+NlAXcrhkYA+8pO0mLkia8UYcGbNi7b8xhDY+7ucW
soR08UHe4bOZsqXXLEG0Du9ObcNk5ozTXgQteN3E5T679BzG6VtumUj3Hl8MfYHSvvUnVi4ZHjUt
2YLml2SlqTJY1JxaIJKTBazwSqGVu95S/oiehvs6i9YnhFEUudsiReXaTq+9zg9zZr+67jAB+V8c
pQeo9tvLakc0Et1rWg3yeY0WVcEI9ThIR7oy5fy1a7aW62vk+AynNW4fNn36UuxJVYimo9U1Atd1
EKOtnCrfqaCMOj2+/AUNV4/txUcMDbykfUYhAn1JvN2BaQdv75ea8y8Jcl0gP+SoW7WlPsBc8IEI
Oj8XxC/0N81ZyVFuiuN2Cl+6Rh/hzFSnMnLewpDSvjt7pfYRs9+v6rdkLdiuOmAYZhwXAtSs+Gkw
nukKV+SnMbjHceniMpxoRNIB4lWXvihuHK+9uzRuKSURGKVkYAN/VtUWoK1iZa/hJXM/AFIZuZS0
jCGTn+qA2un+ZA7dGWnoBzVhYVrobJkD+XytiPloTUeQtUqwaM1+6HNz0KMZoV7EhcT+mzFwj6Hi
Y16AhvE9ST/k0LBK8PMlI+2q6Mf325C+eKzT1ahaaOTgoB6Dbfozy2AKnu0zg+z3xTDTPfBeGj4o
irg5CY4zW+P9Jz2zGJYhBkLpQ0YFQlv7DdqMk73wK/73NodpEd78wbq1VRMbeun7zmDg9ala/ZFR
HJm9fo9QtggbsIvV1zqHIR3FrWKWUtpmf7wHLF12mPDaqvsYEmr3K8FIbzuvj6G23vRGY7kVDZe0
6n1QwcAWKDZ+ZcCaUw/S3OBKpY9GxeScITRmselFT+9GVklHi9z44P4v/sC3sAoiaTcnd8Z+820R
F1jV6p1KGnmVb9moiitdTunkbeQLcBe5MTHa3Qmm+d0yOqajxGPJn4eO2nUSPjXmGMNwCsq80Q7R
/F5Aq0+2MD3Z8lixq/aclM/GVV/0SW29tRUI7o7LVi6Hzcddf2/aOzoZpfNtxfOfPzjDrk59jonz
FoysM9wJjapsvPp9NIao5acN2zNsjnejvZzFI32OoK6LMEio+P7eAtXqbDus2HlEyOgsBwXMyyK/
D8YV/uxhJnfJDDeGUQVwPQzVBWI8/1XAW931llnk9j83WN6VcSN/QHpYxsRPDNvi6Rjo3/ocHb5P
/fFY4Ul60c74nC9Uu+zM0HwLs0vrqJOOGtl3+DP8RLvXteBUE2tyD9PZ5OFub9tskhSNvDe8d5WR
fluIIxRt2Zakvxupnyn5YdyxAfu90o4KnWzC8afYAZH5M7mxpkRaUOsL9WeVE+u6gk4dS2DhPNm3
ou/99ZSetMM/Hctn66jTivIyJq+6RARXQN5AcwE80jsYCV5Dgip2H1D4Qdhlm55gYc7tHJ05cTZu
UD21DPQ3eFo64+y8voR5eJxbk5R/+OQ59XFY+2iAt4v25u+Q3EUgsfx2PLOcdMaBlPS8aHgqNvHD
0rQVssIl5B5M+wuiRE9ypi/CbDVQXYRIK91+VQa2xV5MXDS8xzxLgzKzYXc6fd6svGyMK6NYd1oc
38MgWvg09XpU1T0HGdt29RIRxzTn1wAczHRS4WVrdLZlsBtW6Eth41oQ9bmKZ5CtEJtVstLQMTv4
F7k8GkfORvJECy8VPFVk82FKGZYtzL0uKwutY5ExLnEBtV5mhEaFTQ882BVEvc4gC8qrs7/DolA4
WOWKG8XPi4bEeFmmmg+hvtqXV01uMLGzrHC7FxT4nyoMxfkFyRRxBPPw3FKT/hdTmDSvizUFmhRL
dNbUE/2oK6t4+ChleumeNgLZ9abIaT8g6JArmomJQfdOgLWH6ezLGCC/uAWK7hc75nXmyhop8g5r
OzINVRBVuNJj4tcEnW+oHBviiWX3P4991RpyMxgLzEDwtwxKKBM5drfmmH1SUssUTVn3jKn1CDQg
YMpxyGSgWAL46CIgU0PRbIVdmujzAluHGd2r/Cw+AKV5WgbntWlEFrm6Yw1Ss7iEFITuEG2b47LD
MdNQ+QJBy558tENKtRDSXzffuDiWrSzcA3sx46UPWCtpS76kQwbi5F8rv42pt65+pgWn+Zar1jvd
ns0lvuTEBFHrB/ut7yslXVwmH8/7uDDiBy8g0Lm+pXs0Lij7aFlx4Tvnd//lRII5+GxPRIA6a4S3
lk2+I7ifTeCHfSUazGS7Dd7/KLy8Cmc7/9e0HSFw3FowBNc/rTKclHaMoByB5UtO9oKymKfzOaE7
/PE+LugjwWEAVA/5EHhIHJGugp1wEHpd++FuXVRoZBSN1X3OnKtTvd4dzuYgkWUqLasAYCTME0dj
tOMwoVgl0U8LO736LXpVtdHVMahFFkkyTVmFM/ZsBUV5AG4HZ57nn8WcdK7MXTloMVaOu1HJ7d1K
0IkXZ+P+FlEOL3EEFHLv+7S1hMTg2ZE6Y5eUTL5tSEEu6CfDxFBiobdUQTmZxLYMdUWIIdugr8Iq
Lkf1VJfxxWnCohaHwJbO4JwkmoKPh+h7hitYu+VhprckPtaPY0Ovq6HYOw9KkMuloIXbSHZxfzVF
06fzh9QIo9Jg0qGE3wqr3gWosCygkSxn1P1LeTssh1LbZCABUYXz5Xm5k95SOLGvdQ49od2ew5Wy
E1KLFEZ3wfbiDdi9qK7F1sapzMxO8ZoggLQScIcLerSPyi8W3Uo3GFDdxL8TgPQE2uVOaMSVtq2v
3txAOjXIzqjqy4fybXv05Qj5VLR/aFtZtAuBJramQoIOiR3U0QGOBtvWkYWOicvjSNeLOC1gzmIz
lHIPN/aBztvqWuJltcpwOKVWgYNjkyz3LVR270684/RhegTzylnbVZUSwtTEKDzVv6YIUZ9uCtxn
Avh5nkWV5u0jIcJkBAv2HBeH0VTZWl4DhUjGQKns55+60txmTnWOPklcakkit5Mc3pNbrsYYHP7b
3j/QE9eVqMaN/VrJ8Bje8Jb/UX3omk9tLXGgj11fwafUFhnHGbAL5GfnM9Tp/M+ibMJ7SpDwUe+D
TSBzPcJr0LXYcf0aGqgg6hsYv+jkyKRK4hHfS/aBZIshIiMuevm9p2FPMQinyJCERGVft2G1YrU8
fwhrBsHhRH+vXRHi6C2FCN8KRSIhZqULZvfjaudNfaGdN3xsOfaf8xIeHF4bL8v8Cp7PpiJvLayD
dfJGfjadM+4d6Sfypke75HPCXsAzOBA8RoD19zDo0ih69fiS1ryb0w8zNXU0Kv80HZae5F/nsimB
hAUeJcXsfZj/+Uft1ZU8Td8lxUBNxniggvEghLYQ/cA3Qu0vZlU66sxIH5p1da3sirFhJ7eFoqdQ
HprbankEnAisjumupHFW6iydkxp5jR0bTgbk4oyiGZE7MJji0QDh2s+OJWP9we3d7+M0GphWUfMi
BeQ4mY1yK5z8YZG2Xj9b4VZJD7Wf3UZrZh7NqoDlQxe7WpGMysMB/Go2uGVyzQa6PFTppvQh781F
HeB9LCWvDHsz+l2EwhNExp2i1kUmaqodH04FeMF5ISZORN+kiHfrjw/BepR1VyzdV3lEkY2DKz2S
N//3xWy87MeJ/g7VrGoHcgSV3nLrBqgUyqLn+c9QRQL+avEcGrYotrFgRSPYy+foXok9RIa7LGUp
F/HFyp8kpxedbBrrGh3WhrAnMSsnqq/ISNBCjV4snwE19miKrk3l++844cXcoIlt2GGnmQzGxpfg
BbyTmsvOXNNNfCEjv2PSenzVa3VPeN7S+JGjBz90hjHAU3cHl0dR8z6SX7EkwCLLAs9GW1Apkcp9
3Ln3H10N0j26QR25K4TNZqIUBz489e5mcdfy0ham1lsKQA+9GdfdZiVvxUPwIKZKw8S8Q47dgegM
3wqXoZ9l2cWaJ0fvTQkYvUfxpDT+PZaGhtSb/UuhdIrnd/HNveE56yKJieW56mn0j/yxzkG6UlRD
RVKiWLFrg0/Q8FPtOLQu1oRrrWYjGJ2hYRjJMCoEh7W+0nSHzAhAVrwqgzvWdNEVET3lSFdzt8Cg
oi5kBzgxWDtrXQTw9lEhYOP9sGyaaTcLM1nmV8rp9jOaZGTEtur1rZab2znQ8cE070NT5PM37vUb
BTHgghAtEC6uTIB/Xe0vWVkzTAzIGPcJXsu04vAhGehoBA1Lxxa1sYS+iX7buuGS7T4nFX/DWd6W
aKpQIgGY8nPAOfoPAWNK2oWCxMMiM4v3XS45rNiOZqzhNoG5NXR3vD1uMDQssmZltw6yZ5kiM3ZX
/8G0Cz37XtH8VYLCceAVzaCFZ3fil09D3EL0BM2pKtQh53mSDyUx3Ws/RFryG5V6r3QevnyejZw6
AMBgmqUZLNgn07SINIDxSnmlVoM28HMGxz9wBFuiMqZSYxJ5Kc2H95+580Kndc3ikqJdyhDvPY2g
h5qIiIoB214cPE03TntQxCHcVGtWhk84J0u62WwaDB9EcrFgSXOS+RzeZVpcBJO99V+5/y6+guQK
rT9A85STAyYts8vU7qjKHrCKGI7GRKN8K7zdtm7mls960vR6aAox0cpo2bLzLPS+89/QcK3N8dOH
258Ajf+b42pO7FzLhzrDGBWBcTnjYkJKGIWRTEudZdJrGWxOmrjIhxWNRPYG+kpyp40Vh9bc7hj0
tHnC+q1XomttAj7rEp9By3a1BVgdmlzsqa+u4YRMG5rJOgXG8mWI+TBw+ilG3PxKm90je6yHLYeF
d2StudFayH/ZMDEnUziJrujzXMZKOkTCEld5wlrl8Ag0S9YJGJP959t7QhHt//54iH0w5Pf9qOSI
CHCs/uyn6E9ZpA+las4mZmJSkEItqI9hbt2W3kXI05y7/CpZFROW1WBATMQj1EX2Qzmz51P70u6F
un+VKbpzJJKRyPsq9OIP/ia2tUBLyKTwYVDx2H5J4bS+Whe7q7uhT7rbWYEAsuNYyVwgHtsIOT/k
wYjAQbRX6N1ULQdcE2lHQWj7m5Euc9PLGg389I9X4ewlHcbqf5lt5R3Vd99b0trASY5F1ycFiCGA
/hWI44zAl1DG/rUz86zZip4WKchLdm213VOSffiD+D9SgAffNncRbWQoyU3WCtj1Kwh9eTKqXz3S
AZf3W0V0tsl5Vq0KznCrsh4NXVCF/9Xdiaaaj/Z/VfSyI0+13r4x3TnW8HaAwo62XSjCUE6I4VMh
o2fxq7qimxDfwigi+2NSEBOuZH4LwO+sqtvifExQCG+w8mEnupR9qyHrY+HCdm454d1pc+kwm7Yn
1Nd6Q0SOs6AlOaTV9RMeJhByQXjB/m8gbkNECOhz3ZsK17z2KKou3rTcCca/bXD5o3EEURxWzoie
cQrPBPZelfYJ0aGIwuh+mJWgtz9UQJT9HLdbW1K0U4rNXOSZ1Um59pfpuQq2vPUUYb7aDt4V04N+
iXArI9pnlC6/XYSOS1sXepFTdf/TZNxuTB5BP/B0AF7A5u/cN6jf30JqzDqQQ0Ufnvw+umsv/3Rn
HLoEkz1LTc4uIWzM5Ez7WtrY2Xjdb+q8blExGbaKbNmNOaU6G9J3A7N5VcQgTB7H+WIaRzkEm4At
OwtNSEWrWUtvBv4aXB+2T+2KAp/OGtd6YTBeilEXw++7xQHOZo1eiHU+dy5AunQqtmbpe6LFYQq0
qcZABdoP6aGaA/Hv9l9X61czoE8EpurRU/DhrVeAmyYWI8QY3txJFLX9LLxSRT1Ob0NXHr6PwJKO
51OK9tMWpCILkvf4HCQstzwD5DXiMaFDQb4I4FYb68hWh77UAR87gWoPhsUT/eJWRnQYzIq9FrhL
XWp5pg7XPfHdGtYnqcWdIhNkTkm6yiS3HRJvNsHV+GC3KB1tZvDcGHHQb6Ut8epE+/xSO95IgjQu
vyMxKtyaJiSxLOVWKpJTurcsAEKh4AxN4Z6a2t1ZI0ZXSQRNU2VTSpbgaxIrxo1ext4KRSDB5i90
1rTPnvliuz2qWdtyjTeEBBr/hgBDQeo/2gX9dutjTpmdRUzvfiGpbahDuReyKSU0f7c6a2VKTxkU
GjNDSmmKfs7YlMHHM1V0VKz2Xm+K7S4BdS7PLc9ToG8+JYaOybYK9cwW50hTn4ljIMQbmoIWqrt+
pZ+NF1uD/mfHoM6qpTz3NmaR4RlSMhtafonF8O+DBSoZcWw7/0Q8oOv9DdD9myTr7cyaziKNUGZH
1v6KWjMC7rFa6/ynBgB+XYGyulrs3fjoBASBBsOwglYFcpznEsrXNz+MFQlzy/108xP22FPKsC3f
fFwOfHPR4zOFyhqFlLGmJACzvtMR3257HMzTvtS1VNLQ2C6Gl9BqEO4Oi53xxsFe8EBJbal3HUQg
XqSwo2s5Yl0TRMNvx5ZeWWAfWvYngYGrCORnTjJrSbPbo7OC4lbZFgIymYt+i2tYeJ+depxj1D0p
4dpE6Xeh11NMh0IRdbv0LTMnnHphbNbIDhmCjGqzzsqwtxm8pcOhsLCLTZ2DJraelxTxJ6ueiT8w
HNnTkrC4RmV/ODqDUCwyimizZ4eRG1rQBD9Fd2No72syBrjJ3Ig0DVuIyK2DyZlVOrFJFTQF05pj
X0Nrzt1uFzsusJfjFsuEoAosNbTWhbjiMGdDgFFH5nc2bMV/u46Yl3inul2rgC3RYWXgqBDOtxZR
y7quCy70mMYgfKxsggVv7UwOCdu+f+iUbNz53kTcBT8uVbX8tHkldDD2bZ9ELRU8X6JSRX1ugMKx
pRYuTsUN6q8NNtVOilkBldjONsF0xt/ealuRO2kZI9ylTYt474KWIHk15fXDNr2y+0eLhDEYRm9V
vteBvg6S5clsL3QyWAsY/Pg8ZS6d0E0LPwoyoAm9lIp231kM89QNJ0cNIwdLJ/1X/+6mlzN383Ih
OeQKiKljNgfFUHqu1wGFZIxqxKUEs9Kpl0Z+mP/YRvqPSoQSG2zPwun/FfK1rrJoP00Nhrutc2dH
2+4vimKnh0byER12d8huJ5QrcxVbIYFiKRMZC9whPADxLZKe8jl2an03as0/kwb/Eni2MjXSw2M2
7CTodHnBPDLmgzozIIkqDw3sPjE7rVmg+ukPvdXBWpbxpcE4cQwcWjKFOtd8znrEYGb8v+ZOf41U
jbuMYI/ms/W+3E2oBY4hOLHgIFVNItQ66LuyaQMIrtAjL6gQA48BCCkqrJAsCC6ZQ/CHZbnbqxXU
knXUi6sn+8v4VRiZ3qdhTqPD5EADdrMClqQmuM5TYS38oghS57jPdbPp41hOYKFwYB9/8j3kWZsC
qvWRyi3JXq0supp6WjIi74gml2+6YSpINM0/JjbX1484HdLSTW3RmR16+vtaIB5+EVZJU4oHLL+/
ppJMHFtsIx4dQZYqsBEkNLFbNhQBTzVEUJ4blkJJPoaXmY9h2gTNNwL9EVbzggy/wM2WdJG1oIky
YFo1MMKgNwqnAMY0U2crOg23cx/LlsSFllCuSyfF7gTtuAZ4UE57mJ9bVwIoWTyxvVP4mSgYPh4F
Cy/Oz5bZ+IlNH57JCJiadNC2XCT/NCizgat5y5WTmsQfjy3z5KBnOQGHPbe0tXa4c7+96KGqPePv
N79Bo/Arn5eNHLWbap2pIBEXFMf96LR9WQI82dbAaYUT0TGWVhdAnKhIUV8ZA54mOAs/4jLD3xER
iP55lEZBlQwcjqUlvu6ywgpgGSrARixGTCUfQc/Mla5216OSxYcVuUswIZGrHqAeep1y8m0V/CbV
Fvy3gLI2PxwSV/LS+XyJ6jUCgBH6rL0AkUdn4LWgbapA6vIuQKIZZkorAd/OUiutKBRsrX98UYUt
E09OlYtoQ63ZYW/QrD1g8JF0iTBLyLjEm42TrTsq3fMCFsTR/aWGqR8k1w2kRbL50u01HkPlKxPx
04/Lr9uu1tgZbDUNphuVC6M8wjimszxfDSOQ58+i6ihVkYxqTdcNkt1ewFYR+ZLL+dT4e6e4h2m9
dH53d48dq1rhJlFak4beH1TO2V7ciI6tmKHLIZ8MJP6+lIWK3j2hPY1dSfxVJwVVvI/CyxHObrd/
QRTcItzGehBPN/OBNiorty0DhBp+bmWrMN4XAPmagu6kDeFI5XIQmt3Jvaulu4ROjtCNGuV6Kf0u
KWqmRQ3uhLJMYPucRiBiTLywaFr9Z+ZgKzX7t6+LbsvMBA1s0vwUSL1S92OUlJVmkrq1uP8U9Wsi
3t6/PME1uXcqYXvvRTE9dR7KToVuKOjgKZwmzWXBAkeMJZU7zn0cx3dNHLIBP9TJuXT0n0Qfg+D9
lodLUTSh7VORbBAzVemL+zcHICaiek6mtosVmSgh8N/vBB8qd4HgoFgIaMMuWiCXcSF9K3cNjlwx
hz5jYfSyku+xjYMovT65RE74UD9ETHzj/0jeH9AaZMUAlA0clkexuDI7kaHEFkX+Q+uumZ/G9kgf
tcmRLh3aJvmf7ez5P2+eSubpuC+ZHMdibVy9Ig4yNpm/DpKh+2sUpY1qn1n3Gx9JNFrCq0QvLqcr
NdFMBbC8vEuMGeINssO6SugEsDdzvHEmzdXMgDT44hb+VEb8S5qGSba7TWnqGIU+Gsuzj6TFh7vB
NSLuKD3FlCOI+jxIwnxfCgQyvKBKTFsgs4lUj37cMjo9u4TYz1oOAaAZFvvz4vf4r50wm34OZsb/
WBwc+0ncXW30aU9sBKQmkHPH0+CZ1A7RcTQDoKf32AgoMYcVhhbAfOCy2/8VP/zkkiWS/iRzCmPP
fyqAHqJFqtEr5+D4/0ztsWCAM0gs/Nw2JicrWmIEL9VZUs+oRk9mzJObcyvxh4XJJ6o2lgsB65TD
PNsAedm5uk2bA4IQAQrDR4TER2oBUF4qLmx/lSc7d/lxotoTja48BmwRHpIFnt+AxMmb8wvcnbId
QsuEZqnpxk31+BHVFFbApSNb/xtrzZV1/dREKSLNaY6SusNSQcbAqtCPy1/gZH/ISF8AO6ekvjlM
CDAwnTlH68wmqeENivRgvWOBYtoKe+fzis73dv4UCyBjbH1MbDPxIWmU6DlhoIa5I/B0FfU5WGma
0Q5MI/CYEL/3LO/cEJKHcNsOjTu4NP+LK5UglXa1PpXnVQlpR4KgoP8GAUvFU461o0lqJJMAnowc
/5r8nqLC7edQFs5fy5iuYVVY+7R1ZoSjGvezKgD/UsxzSxFRi3IqwhpLyt/SQCKxn4mVjfj5waVb
3AvQAuN+GsBX204ysWxHL8HZwyj7MwxEplcVd0IWUoCuA8JXUzXBHRWapbfjrifLTAHnkPdkH0PD
L3HrChEmn7w2NgnS1xxH3qNmiCWedxlKWmfO1F0+BnsZSA1DZIuQSRI41lsJ1F2g4tLLukkEvxDP
3xJapHPy9bd9Yoom8QZsX/uIraZvt8pJm6O6HQfimwBP8ozEa/GWpQ0ey5JfcMS0fOKTY8fy+vLN
eLRewoHlCIFG7v79/ACV5Otk3IlwpTzeL50lrwNJtRion+UmlwqawCQ6I6MHFVONQ5k8Jjb2cpj0
YsKKjoD7DIvRfrlVXQukI8wKLucI3kS5HgMsSEmVCjbrLsoZq1O6UOxFtnsjS9XH8QUgvIQNp9O6
MKp6h8kHtZ0G5EwMWf77GcMbYAyNoxDIkP1U7vR5GonIxhmvp1PVwOLL16LB0LiJVUXbXz+F2yRk
LIRNa4cdToHumMF479iJyWy6MvE96InP7RPWA971S4XY94XjQRO4W+X3WRHznUgkY1eg5qmFRW+0
eujeB13Ixh97EL+3qTjuy+e3j4Mc3WvAlPEmPZSWgQRe20EoK3y7oaeYv0zA+pVYMzfIHxmNf4lq
BKyANxyLZiyOKzqZ+BhwqVR2QycKl5KpcqxiSyXflf+sY/vZgKWBX85p8d+0zstmknbkF/vjP/1Q
tXbFQyhD4blwFRgmHZm9mocA4MmrYRsTJVf7zmUnDEvsx7RVXylXc+0WfKP+XOOeWYgqkWh8wYI3
Rv871uAsovnEaAn4KMD0nMBPtc07uQV6PbKvsiZVtZOftbbepsUp5e4rSSXQn35Lab6kIwDAuzti
3D5asOQy8n90iPB0lATK9JcJACjdxQJr76yH5goal6VRhyBge52D9R6H8oZCsRfKh8k9txqnYekt
2GgYQZYR4uxIVX4ZK05KIp2FxTDuNqT/Isb9VEp6CB4OwKk1TF5BbOovFLJlIyVTdhiXNP7pFsSV
RxibCnwXlVMy4BniyJgC472E2V7MKhIeef7FuyZvy7mPUqlYPuy9s6xRr9QkEwJNxhMhPNTup4qr
EIFa+92CgHofmD2QuCMv2BLIBttnmJF9/LVGnWENuiKAeZHR8sNYytPhwTCuaIIJpjeQvJZ2pvjM
e+AdiGbrAh9XwfUZNbDBuV1Bbhb8FdyDm7LHwnnScZ/0pYlV2oWzqlOeAveF4NqzFw1EmPGkZpTK
+yunY2AmFbBPEqKZj7rUxGn687B2h3H/sihzq0bCq8FkQCoQUKgfvj8EUm6/SP61Dg9tMrqDqH0x
MDZFiwR5+ULbl2IuB10fappit6sc/+E5+qnFDTt3bAiEDQAzCizoeuZDbwXENlFdQoTU0oVfnX8X
5F0rS947f23KFOptyLx+U8dNas8okd0nikXhAYsCg8qCFIHQ/udWIGnLwZhH2GaIfY12tzsqE03I
7JTNirSiBh3Bi4zGd786jOl9u1pJzNKygzgE+EDDMBYyqh5x9TRSim7m/gesreotg1EgZgvK4OIl
imwICQ+WBMpgKXfPyjAsR4+VbKcYvkpRtDBGIV/GK1O0Js1GtyhaG97yWHD8FnfjLlhw+wm7964k
QJzV2JJ2YQjMYB3xd4YRI0l1kiB2a5r4UjNEn+mFyN3We9UFczQ9pEJEJgOXxybuGlnJu0lCkjXl
poIA0eOnhHjWkG2mTw2k4CUWdZ35pOeOFvVrUXndCcuvCgsCPHqBWZmadA/z2yHKEq/g9GDokZ2n
2L49vRhENdVbWKJa6sHE2dIY6WZvB6KRqJJ+NqEav25Vi4KtFqHHpAdQsvLqFBVQirwuZZ1/m0eX
BHrheKqEUoeOSncO89ZWuzCqjKbFpBqXI0abkCvUZbBkRzDUSm+hFwxzvX4RBDhaxfPWOThCmeOb
5o4MHVN/RYBIFoXx7e6CYz2ZlO3GmY5ygNvxZJQFgM+2kGWaASbG7MKxX89piZp5pniHmvLuZxh7
Y4xFcUOvbzfS1E+1XGdpBfhldAzhTkYlKN6eyR+s10MXbih3LsWfAYPJbX4U5Zq8lPmPtD+2vVbV
F4rD2UHjdYEagjG2b0i6ApsQgQH67LAcXBy92f7vW/AYtgk7EAIHrdPVt42aahfgyZVLc5GYpKqx
yltPgCTF8+WzTNiv12dqR6qrPzCdfFrRc0Vxet4J4Jg7oWgMRyDj8IKC/J3ykvFBCHOVn9ANdewC
mfeWtYo2WyjKlri+0WYXDY6MqOB1MtDuqSY4lib6MscXSiviSGKlFgUd5NTJuIXgzyYls800oxDH
HsUobEIIZhWj8AZxF4TAtb9UzeaVm/jPCoGdvlgqBC9Ut15JD9li2krPjZh5JICCH7t21Sv5XqaJ
DDhB6cRIXUnbqtGMrj7VqP/7PqM3jgir8VJuDVRHp8Y04j3lAcguybGLIkD9HZ5i2KIO5pXejjbK
LnrvfFucEskGyf7DFyaKFQ+GHNRpwZCylnX/ngKP/JHiucaJhMM3OokdDn4HdkbEHCqgUkZUAkPO
A98+IZ6rVLYzQVaygia0EvMEaCG3Wb8c2n1vW36L0p3Voh4FIQJ7p/p0KuwYU1hQJDhNrT7lmWL0
ml/ULXTDp7aldI5Ik+Hw8bpqsmCMZPY6iqJ0ZVUPUl3d2ZtYAlNP5j13hyXX/hELsvXjnnqix630
ZGjE7O+HWTfm9k95N/AHs+R56itKF4d21jCm64oH42OsKte+Kvsq2a0zp45bXPvjyuQ6ZgVM1U8X
Mmdb4Y7VKkI2ze2YuLSv7vL/9aHQwwGFLNxygx0fu3ytcbILJUBtGXppR+FltsMCt5pnEV/LLGpT
Mc/KR1cSgaJC52elduM6uHqxGewSbVQoTNlOSzm+q1MEuvIKAysomG4pnjnt7y8wctWMaq+a9NUr
YZ3HpGiNvLrR7u5v3tG7eHlc7+okGUGnYzWEIMKowh991Noujrp6C9ex0mPdBuS3KBuHZxPv5vJ5
OqbLTzt+j+1mSeiqAYAwKDq8hTOXtUk9P10fTkzVa9twOlks/pRkOUdJKa2oOFitxV389/NhafE2
LoEPYJ8ZX86jRup0S0TAGOG8JKqAjembOnBHGxRPmxgklk+6luFYU7Y8HSL+GzWpIn33zd/ihNL7
tu42jFzTNUUBtBiaNTTTS4CKiwxuv8X243UfC3HHY3ci8m/wI003TLvkG7VLGmM/5CGDcm0d5gvt
mSy/caEblo6wifCE2YxyQhAXkIPfHFTYjPxM31Sps0Lh+MPFUlrpluKVP41oMYXTnQ8D0XdLFZN0
dWwEVg8PHeaaogSwkqPqcR/JyyTtXR/bqWxKTqq802ZLbPA72xeNwg7uGLjvZsNTWNMAOoYHV8Qt
Ij4eM6kaDBnXZlrBf544pt6JX98ofN+bp2iDUIPr2BmbPgK2lcH2R4QcbG1XXPtEOi6rOCK02ULh
2N3OAuBRvNjRjuQqmgiBEezAIYRZ51eUdbeT5nu4tTwOiSVC4qM2NftxChtKFoKwlS0KNohvZLxr
z3nhH9Vpf1X4/sT+THEpzyJ7abNm8Z9b3vgjVXoUKMtbtSlL1bMO5qpLqwQ7aXO1qBibQ1apvy1S
MMe3iXB6DU472x0tVr3ozFhEB6dssmfxwyeq/WSZHPdBqFdrdu0XeEjTCOCahDM9g+UHCQXsrENN
FRBPlwmRzi31m0a0McqiHuUiH6W452fpRKsZdIWDwx7k0XMEe8gdKST9DD50T0wgDpGrTgTQ3/RU
aqC+B7/l2UD6fClEb/0oyyXBu8dEwzLaio7PCsYXaDEQ1i8hcBv1i3oUnPZOipOTdFs0Ws1yngua
DiaZ3+1/4O7Bn02FoNmQV0TTEB6EJJ/+etaPAByOfQkUtLbx+1lI8zfk2RfPzFstqTWzPeNS8gAu
8ZYk17XCzJVrBoQEnpAVWS4xGC9BSFgkD4Fi8ChBrmssVIL/+JXsZ0GCW9Cz0Qm6yjJE6IKqhBhL
N7QM1pJ41keNhKJVjcUoJeg7nz8AUiyhVi6rVvBl0TlWkd0suL9zp8R0LACx2dInZmC9zXZWL2y8
j6erA0LH0fSlUsUgvi3GqhTMSRKwNfCJdaVx2uJkSvJgbi+caDzah/r6wWa2jmznvftQ5lTMin74
6LlvxcnBlHrkZ45Ii6kWQvafKBQWCBqX795tvM3HMOjJmWSuMyxQ/0hdsS5DX1aR87Vblee72DW+
xLdy6SzgQgbipl0O+H12tBj5ZcMC3nw9jOVQh2xT8/2s6uL7Mhuhs05/FdycaxS3+gjZOlmN9btL
YGNvdWO/UJOyFooB+7t60h4WLU1qRJ9dBryFK97xwWByB2sa1x9DGbwxl9ThL5iWODL0qHuJPEZ2
j32Ueo+efkKNgbZLKrrxM7ame9Geed4bo1uTm6u2vCSGg1VcajXZqDB/SOZQMqgQ3Jj+di5Z1+st
53y/H7xRWmohLUZp4jekB4N9k6XxjhBXZXuDNynIPCrReQ5FzrwGGGcTnIEfs6r4Mmh8u+7lHtYM
2k1HMI5DYfblRdtpbzERnAtpR5d9IUZ+kRDJLbPKF1BAz7cQq90d2IUM3s8r6+8a1RhPsx1hZOhY
KkKZl/tZO4cdn6Mtr5unns00QzVM1IsgiSdmZdTlm9J0x0wh04chsxK9AICd0BDAc2MdIKgKLYUA
Dt80qPUwYsS1UIMKr+DQ7IuWVrZa3XM/0zmNx9fb0YKPzZDHhhC+ec7609THPKRQTHgJ7BWSIoSR
o8J2vXWcTwvDDnjpjaU5QFHAd007zKVnwdwffvVu9eaxHkJwh0rTedZVjaWThDYj5k9jd4ZRvbX0
YZaDkHj60GGWKGe73SCNaCPCHNBQDj7RYXwZ/YGx5ZKITI0pz1JLaIbCdqG+vbHDXkTzBHaPFxLr
FxmyxezHh6ht+7NKEiJLHK40IXyAEue0rlt/bPT7Q0pbBfHjshOqlOxuiHSMSLkDcLF9aMcPhXVZ
XHoHtfQpan55YNY+QE+xsA9QrS4GnEX3H8Bmh2FzRRQHf3l+Oxu6Hf44nLEy6BSXygSdiqkZeqnF
xbIK+4DEWmL4OAtHQp+rozGe20PtPiyADhLBJf0A63VSk+VPfknAx5TH6zjC5CiVYW0eDI0N2W31
NxRQ80+C1oBw6W4FAeg36rt8dpJxiwfOw5c398PvJC2HDxojc0M0v2puncDLHql8sBl3GgUI5d7I
W/rfs40MeREPEspuuUQ/dz56gHShGpNjba7kzB0ivGcM3mkY9r+H7GbtJ/Wa66PjEzrtaN2ilfVA
UcMJ6KZpc5cqMRC30bQmqx37VK7o97/zy/TnA2xRxl224qXvSGfMnB29JqQZFud4Dfacav17VtH7
4tEyR1taTubCqGTPq5DixHreWzZksPxwuOgVRED6XDLE3r7gOqvJmhI2uNc+dxYWsUMisTz05Man
U2Fw0frPrzpTJXDnbgjgsbOd0KD7AgjGRywSK1PwzQVlR7Whq19Arr8c1V0K4Z2BuQlLZG6MR+4j
HO6k5jdh+zVjHI+Rpwpqal7PZqifqOdPG79asf5w0W+Mr5gE2MFWwrNgGQ81mD0frn1YvyO4jh8Z
ZABh4f8dxpbznpzQ7GRzWw3c4C06qB7MXTc3+CWFk6dIEQNyAjANRzLnULljdhtTTT2QojE2Nr7f
6f/skSMKAe96miTkA9+OT4uyEGnriHq+/hVxpoLc+EMiKjCaIn/q4ftXoHdvo/ozXXHFF3C4vkSR
rlM40+RtJrB0+Zp4mNOJEiyAanXp6AAR4dK54PDKeHbYOiUtl0fb5wVeBW+9kqXlxVeK3V0vZkCY
zh3IiKAQe0JHBcDobofCt82QHC/lDXw+/4V368VgkvN9/Gkozr5EPXqZnDWHBggaqBkqq0Tw/2QZ
4WjR0C8H1IBsfH5D1WvJ5JF2gOrW0Lp5udisayN7aHPjmEDThf2/542vc8u/vezgUTZo+PY6vLNt
w2iDJaLyTVk0Si3hNuAxr3YZKbuPYO9cXyLj3sQRtorQ97dIMVGgO21HFHwDfv/4+jx0gD+oL2xx
EyjOysW1Rt3YSnALY0GEXDRDHM+Wx5IoRhZs2c+AHn4iq8xztUdhdzq71DfjZ26PZBotIq/Lpt9F
Cw7BdKp8wNMR68gZgw/ErYb13O0xNiT7gORc6hWDwD7mE3Sh21j+iA/QsFtk6wYmeTbmemdumtfo
eIb8qKFKHVcel2vUA7GSaDEA0XaTQ0EgUdbg6XrJ+28a2780B50P9iq3IbXIxyomHjbqEpKaeUVS
eRvMhBgxl+jK3DzdmF08l/eHLL/9GKwSIcQjfZBgpZVJOELHlG3gXbySJfWtzu6HDA+SSmHkjW3H
ztkPsYadH/mSC37B6Sxc1hbqK8xqY/uYyXto0o9V6981I2Q3HOupOHOWu4qDCR1C/oscGrBlOqpl
YTUdlOocT5wDcLH25f2C1KoW8ucPa1bYtBrLTa+nHnxzXVHY1G7S6/B2Wx/Xy8Ph5nZ7NbMXXK9l
OjkALdXXiwM0wauuJ7r4iDgfBS+FifhC49z7DxGcbRmBfIBZUcpu77dU3SbaEgJZTw3+6SLY6mQp
g79FXDSTWXAKYK7CjYTeXSrm6PZU0Imjyebxgkc6lT2L6NidPqrN4lsPoxudXiDrEaWjXHH2TEHE
HXoemXW4J75rDbzcXOnwW16tWiTmTEGgRQt3DndFwOeIUT7W19BpHMGRns/6rgiDC1QN/o/xswoK
qPl0QDs2Qx8tuJLhwIRSDQGiE1N6qEUvL2IqyLMiOd6GOYLBRO5L5KPBOSRJU0SyfVsv3SVCqRH9
KqAiJUjmfaWsl2+irrPYcJCIIaqN+SKbaTyu4NcXq+d29hXt5meii8fi4KlBVbprptXctLnLwclN
8No1yGMwyemkjCkkWfhN7e9eTPGobkaWjdbpZ0YNA963BC3ogeaaV3egAJKcumMEB/wVQYfbXlMh
lt4NdVdwKVzNKJXic43S4e27R9RHlk6P5PCHsrTfsRRhElrEU51WqChz7gw3gQB5lBqr6waOJXKk
VA/HrCcKh0t+t6i5kbiAkv5jKp7Ky2oM7JvmFQmQ5/s8+wW7YeX/ChsbCZLqtzY7FzXmDOhb6bGU
PBFcJYDHN+1xDHmkh+JlcRUGhvrdDR0xb60gQr8StHtslldjtT+KffrPqRs3gmN9RgBujXWXVC2E
J0haoFMR8+RnjTgdZ+RoJWYk5/4GjSKPv3urbwGQro3j0Xv+OpVXITAHSwqfOSbNOWbqRGwsGCsx
wsiUTqaDAx2EcDCN2/nifuZ8yeQh3ZtJtml8r1c7gPdZTOhvEFfbPMEtFRb7qyTtICgN6dL6M+Pp
aGepCpS2Ai/UKDXPTrZZRSTZxA/CDnS5ECVEhKfa3+HvHewaeMIUB3TzSco6cpGz6OuJ2Qx4Znlo
/+SgBcibkxA1OW9hSL3KLTWUx/ZxmPAzBVRxr94nIqI4RKDc/y8DIC6Juq7X3RO/lp7jkhagCP1s
5jV8Bq+O1+ydVhz4qJEtyyLpJBFslHm4/qAB04+mpXjgM3Ci9vl0AsBh+xBA+dZ8rqlBIRPDxgUR
ZKu2B/fw8VLOu0G96xLswp9S4aZSpAfsH4pTLDp+NfHO0YjNHHqFNwcsFm6Lyem6rSX6zaubLUAk
nCDwW8eaGFzfII0fvRx7GY4g1X/XvMisj2ZGzZ+k0knPqfCkT2Gifg7b3TKrwOqIxsgxUtzjErUA
faiKd3ZgHIZjXSVcrd9VfFwJQxJ0tpuVLPmOW6tCE01wMEWf+fSFJxqC/3pJYNvtN/dpmq3UCAE2
/AmeqLv+Sk/GiMO70tL+HQ62YbyxG+SKFFU2BzN+EDqP7eEty/Crsryhb72yV191vYpctnK/WYGi
ZRd+TOY3OOqnETJ8/xR9bjm2vOGuEJd+1YKQfzR0bVQPIWaSG/hhmerkgkVLkQHxwXCxE3v3TzRm
Qer3PAv3SRZ/hzD7FA9MHJc5Ele7MkL+WS/C8ArLvlkq2gxNe606JRllfWwuUeOLEsBe8oslfQtf
zPWzbJte4jXo8RdemftBbmUvIG4SGFM8X/c8H2od6pC0D16I0174D/WdVFOkkuF9WF6QBZwRS7XR
K0ToeHD30PHgUYkufi+KfCc7J2OUvqGSUCmHpq/FXzG0aW20w7dS4QvAv4kMGJukaAiRiYA91VPa
RXWHfvovbElMtTEDu2SQ8v0lLKUEqJr42SJABsIQoGRAXqYvqC9fBHtgGt9YX23cijbYlKJlxFtK
bDCCVSoRD0JR5GrSWjPrvb/CJS7qAvqvTAI00P1DMee+aJoLmH3Y1a/YvHt7A0Jj3v/ABmhobFlI
WNAFpv1SY1zrnTwL5eMyUB8dn5ca82u+CzUQ+4nqHEYdaFFWw5r8U1LbWahXOX3uEiLDagh8xwXc
+VUKpOUeQyHC6s6+leo3IOoJoVqLoX4WGhVbvxsuQ6DLd6xMXq/Vw2oxsX7U/WOWKlrKaBOgA2cK
Ne7C1CVGJT5SDNwWjj2znhl108jS2oirXuLXviA2czHoj/3LNVS+Utjva6Bf3Khxq3foiaRZsMzh
ISlZlXu9CWGs9bOjmr/YvLMzrC+8vFmkSmpQ2OfjvDLkqUuo5kYiBVGLFD4Jfnmi6NLyoJqi5UtF
C/SoK0YI8/GL9uKQuCmkAy1Mi2an2P4jXcGGwa/6YEJpJ6zmTwBYPRMJjNCaHP6p6I1c1hcH5peS
ofVSZfzYAc5qX9SCko/UQhih6wFu4wWMYeSHFfXCW/tfCvh6x6H+T68CjWsrwFbtzblFVd+ex7ma
GynUAvC+pfFecjisGL11P/Hhh2sMwRx1t2KhYwMa2y+n+Z8jRfBVwzPMQcIYr255ghlO+b7Zz3ak
7rlxe4Ls8XtBSdzoQuqw1/HGqH/p/eb+LR/Y2KcVfC1CmMy6YFIt9BASY3tfbYsNx+m6LFtEluRi
CvhcAAU79JlQeq89V8agsX/RPxICONtQvhrlcXOvQJLflw2mOjYIZ06ity4KnKNM14+ZirnGEPYk
j6Ew/b2tUKaf3vH+rPZ0mcV7y0Y4KPbleeUM/mkqqMjcZzjdKePqwzCFrebOLjbQdYGVY6UaXPWy
fp/uS4gu6Fo9Z7BJcxMsKXaux6DyOcak+pLyTief3YaOebl7l6YHCo3ZXIALEJHf+OUgiJTqsips
ldKxUfwa3VF8fb153+GBd7xFiAtw9+N6OmnDAH+n+y/PvnPZ1kZzEdXP32joPgbwAE0x+BygE7go
qdKvT1+tXvr00v8XDoAqlu+0M6jIKSP4xHuA9RwmzsegejB5+hBu3bRV8wcfUUAaQ/1ccLueu62u
ivsyDu9ogVFMRsrVLya4Aczxb62nuAcR7UCOLnRVcmOvwnKOQLswQzOxnLLilLPXz3cI/DEwWjCa
a997rnJwq7QqK1sjmws5oEwaa0EbJXK0ILmRXBW4NW0LnXmqk3wZ98hgc9XEFGVXb5KF+WQFqrQR
VNiLVYipy5jyMP0KvjI2JjneKLi2gh/vxeNc0HVxxYbhOhNaHBqMk1IKe81aJIuFcruqH9twJ9NH
X0nfEFNG8eWcz5fvY5xvWm4++Qfd3uAswWK0n61tQfi1t/6K0d2WXJOm46mG8oItKcszsWhSw+En
6vWWArJLe3CRgVBPX6nSev3GzbfmObVEdS6QlFHuvgB5iWHFGF1Yq5QcNsLsJ45mbHkJQoX+H9x8
vVnRS/BJYc6DAA+5a90wS6kXA0LhPXvZ+wSKDUbpgAKTcGfPYCBS12hXItXdqutxoEOAhSvbMWx4
+y5bIIJsfPiFY6I7/ifHVtg1uAVIw+KIP8TWiy5NpombnEZjiEH9B30oxQmoXI0dtmZO6L4eizL+
ecRRg9NWD8W+3JSahw1ilUL5rwgpoXkhzUj9zlCtQ0yJoMC57YCoU3cDkQSYXVlrftlPBR1BEDRU
giMIzz5PNfwuw970F7FzRpLfWev2EgZ1ieezJnj14GQZSBtud/Zvq26Itzo4p4tttBpwnj33JbcE
blQ9Kn7RmRX+2mo54y4P+XrEj4eQTQblfCMOh2OPoJee0nCxMNQZN6NhO+xLIzPKRt3rFiikbHPk
rX13y9JV2sfnGoDX2M7JRmb7qElB0SnLXR0d6rROBsBJHOQFEofg5Neq3Y3e8FzNXLsrgJongLLl
W+ZUdtaQ+sWsIsXD8swIqH4SA0Aor+LJD7uAmBSymvN/kAKIaf562tdW0yb9+pwKi5XzSXzPcynH
5rDmKFKzM1rWAogsdJ7oy/rKlGGEXYJeFr1pYkFtdmPKWgwSOdsGz0tMpMHG0MUBO0MTgI2JRLlg
mDSxsyPDJIhl/gJz89+dRset2sWz2A/8RjKv9xHvaVXZ272ByGFf6rIHRnrz0Z3tcVigouHKGK1c
VwVuFj6w0lj6v+7v8N0dKrb4+GlumGXMzKlL69jOBp+VbeOtTDYyonVZQJz0i3ImTgda7snvyKyB
W0gC4oaun8OEUR8+vzLQYuZq4Qr66HM+Indb1tLQpvu7mX/Ke+StiAGa0DtZOnKPH/+xqeni6rL6
CZ/QPEnI46HlUgmSmrPrNTcv9fuGmY+23xihCgL1axv7EO7hVdIiHJ5Itf4iPDLIpAvYReENs0dT
pDJcIgv+F12Pd0/eLb46X0wU+WtUln0iyQ5Ohkc9zCQyP4LMxnXT7ek7RbHRYpcHyVmJcX49baYH
f574I423bnxOErDb8PXDQ9n+nDUbXmdYs3s0gQpMTQURv9uCk+BwzhQGAOVR3l70Flt7p3b5jJrK
FY3gpbzS/2yyiQw/mnnSYWoyRIDYpu20B9wNZjGr5COaHGdW2smtyVdvVlaTgaUKr0kmaA1gqpjl
pomMrmQ2KqgssDzbuH05I/PS9tTkJrwnHT4TrnWtBU069+f1Khi6q1JQaioA3nWB+JW4J29PfJRB
MxFpL1HV9ipi4iF8xFuxcdyZnK2T5TtDdfQBFziBeUZMUazA/oAPnxtqArCUYcVup7sSHSlfdmuZ
X5kUzMdpw8IOc1Y++87wM8MTlYAFwMhQKLAu9S8ka7yT2Gag0TrYrxLFpbfm44n+Elaauk0+XLTb
vWTDI+KXi6mEg5uAI/+QLMHceaqwuC7IJjyC4BmX8hmRNfhZPBH/niyGKYb+Oxr1HNrv530XR9ud
WCfaPtPKQsQLUEZAlAFX4BJ8eDl+x2yCnxWflEKfBf60PSTuMdnkQstoZNlWnT5FEEzdK2UqPI/C
BezmxqWPAsFDjXFYsGoTbkhlKLbfPiFv0KA4lmhcTFIPoKenpgonuaPY8s9C+V5fZo5ai/z/Dtto
NDItxm95PiOX8YfDsdiS4aZkeRaHf9yZw7yiC34fx7WiE2yMymOfaeWPdrQUlSFTQ9MvuAR0xZvZ
+9QoJxhrvfw7uHusyO5FEbBIpdJ9obuPssQM2IVNScKH07kCzceSM4RQR7HpFwYNvpE8bPihG5Qc
+89eCUk9LswJDYR6YNKTnDofoG3LWOiVWcBjrU/1SpUJ9FvV+UzQ+7D4EWcfCQFQnrrxlx6v79DA
bJRc4XGfWdg2TfMlQy65vqGDy1bsTxFMyeNXPLKkbBBHWtHx6iVhu5d7WW7W9q9IiVc1E+yC/mPP
7ARazQEcpMhsOyWR5D4KFcZbgaRnsO6kM/Tp2e5SYUHjdo7W4slbCPUqTCRGjoL8n3b1Mru3caoL
A3H20PIvKfyENxM4fS0MwRAqUZIdr96xlFdTwAvRLGRgEeZlG7nvY8J4ne3yFDRWy19L/fUeBa+g
vk6224P8ggk7Y+Ga7L7BKVJptWlYlUHICNLTsGOUuN7q6gimG8/vshrKofyLwsyq6Atxq+VPiEXd
fOwKEy/ixwXq24habTJSQNfiRxcpvnj5dpfZvhf73Rz2Mpu5VhHCdN/qQuQbfCt6RBj8g7V+4s38
ZieNr3t+wSBqT4dDrcy6CTgv3RLN8194TnyLjV9icAIATNE4HAU+jE/UTJYQTlCNEv8Rad0TCrkb
GPo9PSa2G5ikiWQiGOiKVDvXQ1X8YLCadNnLcX/09G+buYG9abXlguZJxBLAjgAiKdpkStDJK/wl
mEAgdrIVRASPTX3qW5QMgX2fw3l6aOe8Fr1cIELa4NNF3OyRwUBh3xG0wyoaqoAFqwbGoxYPbxtQ
F5uuUcNj3AK/ZVnS08tledLSio3UEpyuDa5296bGG7D5Tb9vvFK45bEMMdljSfJ4Rkw2scGDDqEP
z7ALXi18DfHY5onJXjMubK/2GUIihb8znZ/gGvX24FBbrtFP2RCkhFenNgjD5O7ct29DTTHnT2HK
w7uGhHDixnDvhT8pF1iAQNDlnfQITxdTsdljtb05i5RZbGLDZQ4pb22qyLYn1/yuJPGJcFN7j8+U
tqvBY90vIDu8/BtZwGSKYElGhFLtezVvqs3uS5eMWwkpz7Z/32PbsJ4JnFZD2R5VkNdeRcTRG4KO
Z2JNFa9xQdzUMwSFFB8PQaaQLr2Cyvo+VZomP+qJy5pEBTKB//zmBxFoQTVmP0dQwnEYYavomj4l
AAHAM7HoXP+FOJGWqw3WmHUQnsACh4SwST3bleffQc0y0dn13YyF2T1VF1MlQ1/t+3EnFOlgdUPo
h6am9k+uYyfuc/jQlCVIYvztKtefqhfRZ9qtH8CY5AvhlYAj9AjZa1Dx6X8O4UKMIW06Z4KKFtoM
yWNrIMtSNmcPgQLdNF5yBUrbCfGeQ8ShWahsmFrCaQ/hti+Srh0bI1dg4oH9dmahmvrXCmHaTjW3
g59Z2UymbIIh1n+GGQBXNK0Lshkj2EnshK0FO3KrZbH/ugXTeEhfx35DqXvgW6FQkCyAM/yQWDg/
MF8mn3TYJqfM/dgQiss9su7IUgYsUNWtT6VZ27lPwsn4Dr61JAI3U2YjFWpJH81WGTolLuLktSXN
01nEMCIXsYrrH50qj/StqJ/iMzy54q9Bvz+C63pcTbMM5pQCqrNRbe9oIArR94ikEbRn5qSb05wX
ZW9ogyvGY+w38zvBpGwxp8G/o3hW/iI2OgzNdNlhcKeApaxrVdsFDzlISHPui0I92hBWOS311SeX
kitw3VKnzR4Hh+33H/fAOoEnDqGfsNPNMvoEZxYpYq8dtJMLIsiyFMMroLixS+2UuvFgSpFSi5Ba
6gFU7xSVOIEAxdYCGLpHud9i3m5cVigGCj5Ez4BV3vvSXDvS355fGdSH7yoAT+DYTT416/hbZ2oq
sUnxzRsEQzHUbEsc8nBMQGihy69EyW01xlnYhIQo3/wK8dzgSJymoXl1CLjEmzRkj8UODVVDYKP4
8vRDmQbo9k08FdyeJUUUJmrux5kyIORHjah9brw4ZHwHzqJdfl6NXKLRvPZxGdWOc65JtQYZBXIE
+TyVbyLV5RMXfHL+vfhr0ctV/xz25Fb7pD4FPLFzeCYLVjPUmtq7wttBL/oz3GQ1FlRwoW/b9r+M
3715MHbJb1qt/m2xYfjvM6v6urfmhtPKUDO9GyGIfkP/2E/Ko+q/GFJGRIkSnU+5h5cY3MD5kuim
6kG/eBmQZUT5aD8SzoeCT4TEPcSNQBB5FUJNyvsyazFSq8mmWCEeIdONI8MHG/uJYISLKG4UgWfs
Mis/A3jGVS2+NW8jvGTNPapPwP9YjNlgmPCr2/4kvj3hP0NrZ5ckdtwuuJOHbLBcgljR53kibkgX
V6cxA6iMiPG1V2t1FKfh00fQVTCV5lbXlEOBytSZWoDyBny4rF0FtzKFQ+55Buo0nvMZ9+pP93KQ
AsZa4wkPP5VmnRFa0cU/dEa0LiCihYvK3GvcN0pCqiX0JzNTeugsPSrB4XqkF9AHv4GdXASQ5eEd
SWrCE3h1vFBsMaV7ax6lUGQBHaqwObE1oKiq8wOGLDJ88mCTGmA9WSXth53cswikpsIuZs9wnsJN
I/r8M0TLGWyDV9v2Lw/1jxuoGk40pHl3CWGiGhgFvU40/dASb1N03w3d1yw5I+iaVlZ/jPWZVOOb
d7EiVmsYWaQ3rDbh7QTUvEDozhWwFJMnb/GKbfmhvxt5LJx1kCdmhQjzSuipPo8PiTVyZKmFze3e
JkSlNTzgdWM9EVA3BOZDE5ated8pQKK4CjEWELTqULSNyJk0sffgSf5s3a2QxTkoE861KL2V8oPX
g+qxfJsdHsg4luuzBu85rp+mrn5PB975vpSnMRxSTU8asQB0yRbK4By8uIfEHvvknGQTvDqDjUAc
3YhLbpgVZNQoiSxjkWogTz2kNQEPsHeBDCr6IfJDHL5l9OP+9TsUT1WGb9mfA/DhAgeGOkYuPCjZ
DLUQqsuvP1H65d6gIfjU6IcWEDjDRhw3cDWqi114tRwL/dA8qpzX5z/Tzl48f6mcvStObhGU0QOt
jTCQEBxAhUejLGgqjfwKxY/26Xvgow5GlV/6RXt1GdCl8jKBEQOszc6HmRVeHJ90TE/0AgJ+7roI
Z3ANtBcwPcBiSmyPmkVscDHqgJRXhWMrteHwLcygacsSJJ+eNhfMjHlWp6+ObS/KLO0UjT9fJMog
BLSmFdgs+JC5nRJkotJZpkSEzcYX9cPvrEBZwWhPFzQd7JtvkYqXCkLLZDv4xATRYQgvWFbQEPai
SabjlsfWPUuBPTkyC29n03kkmJVk9+c9q/2Eq1oovVe6R6JgFlTazB/DYQ1VFq8WDrYWfyLAgmFE
YPQDIRjFrpxaRzTDRxOATRGIzHlxRAzaisj0137QbQhWDYyU4cctaVug1gMoMS/P+7P/VfcgruBh
yxYkw7dBMGqScFA6/PsiA4I/D0EyHB0mA7lAb6CTPXwC9ok5H+wipdj8A5urdE1bLbqfgKP1g5rx
TW+O6SSH0mKeL0SYT2PiQ5Me2xmURaUobXP/nLF9zBJqQ1oOQVUB6SCxczjqs4ViBlf0qWi8Tg+s
NJb5H5S5cFFiZjzMj7UplTNE9pi0Kus6TjKnh9MDNunndgR0SvY5KrgijB2nK02p3xevutnC1usZ
q/+R5xRFEx9iiHHVLL7MjLwhyPCJckykvYazDyDYEEQSakB0+N+tgmm9eZBGWUdp0TfyDo9AcSzO
/y4/E35l2sV/gwsIeH4HXzD4MDHV+wJV3z4cJsIhiDDRlPCF8mp0bRrLNCZVuO5YgskIjxmZHVtf
sFptwc8QmATOHib7KxU9hYA+tiStvyOUeM4wyjs6gx8bIfbWJ0gSvG8S10vPu9RUJG3TVTSIlRd/
hbJ8FQX7d+oKtcDW9TVVcNFhE7ejejzpX6BXgfIj748BGbxWCfpBeOq91f/p7mFm8TxR+yj784X/
kR73ovvr0L9cqBIUW0iRt4ItHFjtq5ReAiUQ4alFWPDo6ud2Utjp2A1bLss6wR2pzeGzaLu5mJEi
mbZD9FmJF+lgHbYJ3KT8ECsYiGzCvmh466K32LWY0+50Nkp0JQtFAObvOU812S0F/VE2y+qN8yNA
GFrwG/xozeqaOpC/yHoN+dzpERcVTDx+QWzmLB3BzG353zTZHLwElCx9YuJsJGXYZZb0gHwQQTap
PlgsVNh872OIRaR3RPg3JNH0RauvKbktepKq5FPjcJfGWGNj8TbEme4AUC/cOCFZ9qm3fuLiz2Qo
tbJbeJ3UyWE4JHTG43DQg5/HfwfTY5wr5tO4tJShOxZf+H7Ctyg6cvCxp6IZDoQY39WhFSuJqf1b
pM3ju0bfAbtwewsHT1gLDQukY1gLpcGxhrOhVbInXOk5/X+tDDJC/O5kA8N28Mg08x9Exi0bFaQj
inORB1R8dZg60No6UCQHMwjkGUOY242sHGW2IP5W2KCoSttx6S9vZf3y1ZW4QNqEhR7nLsOkmI/k
/jtNKpT+4uMGYNi3GvQX2HhMclPtg47qndbBVoBv3FUKMcQgFikqAhZ+lY020/DAoz+WjREHwidB
VtNY7fC809oSzn+/REbPHbe00xzogEGkJMneCU1mrfQpkzEALFSCmJH3o4TPC/MdN6f5zBLlxzdf
719T1r/UpmFyi4HhrMj2Ge9YaSYAPJi5vfCIATMVh3mtr6hA12EDegi4Elyah+W4svv16xmYODEi
BUgcUtqx6hfBtCIWjitGVEp233kWJ6U4lVxrruRBt/+k9jqTE5TSyz159kdoLMix22uJOHKfyfSd
tISAD8/anYox3ZwAwpPhbEaSCK+Nt4zx7u3dD7GNRdTBXa0cl/LDWq94/mfQA+crSMnkAKMbcu2f
zVPj430bcnzUUzX9m70Zf4W4bM4G46SgczTKI20+LYJd1x4vA/3koA8eXG/RgKpB/2vQFSqphNVb
KtSSCQx8d7YxzpVe4dsBR7U3L/Lth0s08QbS+g89mHAUoAWKPeJS0zjjpPeAJEgIXnWxS7XErxcq
I50vUipW6yG9undIoTT1d6h8NRBgNUAANypnpN5WfbbJk5ibfQ0aUQket+olFD9CG2wUG0dCLBF+
uk/qE7RHD4X4vfXYyfWNa0DBU4N/0MYVyfKlPBtgL/JH/8pN2r0572sC0LxJgoHOaaYg8+VMn2k7
qgP2TMNDOXpBVmlzcAnkQKRQQhX7blU52KX8WNF1SBjOs9kiXGhbRMejQYftH2XuIR0yEymjdyHo
NL9IqrumdOq/7SI7AlIWV6lMozZYoXE0ixPNE+Pt7CbJ3U9mVvrDg4cbjTCl4m223hJvZTYFkQXc
zlpucKOdbPiuLcc35EG6KwmLxukjyVnLm1cpGrkWE9iYt64vbZr07zii83g3460Bsqqqnt+Jm3ib
L6w51cAkbpudeVN/TqJWuHk/7nN9nIOl+NrKql6pJc+mJhYid8Y73+tu+F8DP6Pvq5+A3GF36l47
gRcWsgTGT+QaLlZeGslFYJJxe+RDDeoaWSJGrBrnDG3v6E38bZoIMzFi8ckOFgmxkmxdgWEZ+z+s
MmUDT6CwJk419iUQovYldpr2oUG2JzVBQ/DC9OLOs3XKbUY4vyTPWUpNxH3JOWOOYJbovdL/MImF
neX7gvgtr1i9qpdc7xyOtmpIAYd0jvM1vJhw6U+K07V5tO9MK+h/g9JMa9rTrAb15IqckyFhS0+I
jgqgpusKXE1vCZCb9T1/UV9kQBY1SMiwXBHMp8EzfPY2Tkyt0EPhVy9Vyf1wkggzUI5//sAAB18+
yN558vferXiLS/kQN7qn5LAfuEooGEVmDxAoXiy98+EZtXdiDPGSI+mWnXk7J4qkW5ZKrxGvn8aG
OQbeFphvh95hmrfIKox7fw6rJ0cUQAHMsO9VTmE/mrOJ9GWi0S1H81idXOhmaEqor7tZ+J5n1VuI
z5nI36oJyPqthZbGbFAqatSmkPxll0xcO1es56DcpyrWPvMJ+6tTwnqbbaH5AquIOoeEsZA+Pf+U
J4X0LNuvJVPPdTaGRmHiGZ0i9onNwEYMeQCVPgayBlN586nNIDVZHXJu6g0Gb73G2fdul6YxXyVs
iTwRxvUh8cQ8ew0P6+Z8D7FyBG9gGJCjudkFXpPnOghAsMj2ZO2dNg3kr5wIWAb8HSf4T62UwYYv
23SHbEnjOYnpc7hlT2dpUDx1+cOJa+STLtEd2sXU0XrFSVJqXPDSawS+PaoVAYh+UX2I+3e/PypV
Gz7iAxAmYDsmmqB9K2WALw327DpnQTNRDRdsq9nmUjsX9wOm0XRyzPlObQfCtpz/JxEwWJPrO5yN
Cc5L2uvJ2GuswnKo90+ZrDH/ALJKmZlwa3Zzye+5/f/i/Kv4HluWPh/4c6cWA3SsB+JosRjDl4LI
IjI0cMH4Sk+X4Cgl2iSw7hx7XmX8UIF2wGlcP6Vs8MvTkigBa0JlQGivXqmoRow+cEDeccA57kua
zPf2nkqmNOE49lI/cULRQORK0olF0gYpBUuhGbIzgbkLHUyXLW06g2tgTMkMGtKQ6TmOXkqiJC/5
H/+A5bwqbWBD+rScSww8akzO2weDyIOYRV36xruU/P4/VxHkCxTPs0e/YdDTfrnlrp0I2WlIFr+D
khf91Gwvfq1u9xMpGs0JNwy/VdCrQqznjDEUQzZYIUGpXLTbZMmwJUrT+XUb3pb69knOqcFP/IG3
nTcngs/+UhsXelnMOHkKlYxt9W1+MN1B3LTBIeVVUhP395STbTnE1g7Ucl3/knnNsd5U0o1TbEsW
rpR3kpdvlKwP/8BM1viWVMOAmSOEWIlsQcGqsmJxqrvnZVhv61Y5v66Yt2CBwUaP7tTCkT2LZx/R
5EI4sSpwlilwylbExszSxGB9BZYfGBweAvkm7gzMe8/l+6H3E6gPErlPqscDzIXKOdc8OGy2yUOP
lhz7r2KoaW8UzSBGzR0jVrZX9svpHEavERdaydmkWkIl+OgrwmJwWyITNHtDQbIw3lxgazAJ1tkI
1Jv0AqPnL73wgS/+GgjuyxWDmgczNVaAmYyfGTTaYJPhQXef1Tvc4nCvKOv2H6StI2sfXDlwqhYI
ShT4ZgV+oWy4Djx1M2j9QTGaQzlXPzXTIoNYSOlnzmcxtQNK5dWwinFl7pO0dGii3sOrNU7aRert
xOEuLAH6PvmesJUyyNE8fMFPsQRre1JtrRVAW3P+knp+uPSqsmtkDPgZOqmikhTc2hSvkp17hCRT
EP6tMMibl7WM96H9wvIGaFo4ORdN3HOxb043cSVbaJKnLmsxTiYbZgvvnV8B1KUDP2P3CqwTGIx9
RExNjAV/7U+wCj8UEg0Ozp+rCFUTYV4n/v98kmRNElfM9Jvg2DLxzUWdV94ZGH7033lmQnuDlUMz
NGLu75Amofb+fpgpfX8Isuih67TNCySHGDSgTMgbRtavK1oo4t0rHxvqONPrIGRff2LdaBsXWELb
6i0Lwfh9yv1id/MSn4dLH/y0WjYzX2aZIjkGhsfZEPPecIpLwhZpWzhfgoNTGUU2Q32n1n9uVFNp
VyHXVqbCK00U05wPawQ7+CnIZe6MO48LXE1QquDyl3GKAsj/HQY/h53JHM7EJK5DE21H3aaZo3iM
fbAb8dclMU2+HncxrC+FxbxF597iHhHvDNMXL1mTRZIUOrFFCmLFHfz5hPCq+4zUC9WYe69Sl5xQ
ek22V0U72Uuc8RmTvPmbYVZgrOHXF0RuXGkLoIHsgzrSU73wIafNTI8egh8pVPiORNFmfiHUp8tk
Js9TxG7q0QJvtUzr7zPr4Gv9BIRr7Vs+zIBCyTInmb+Mt2eN35SFj/uKSY8T7fqYYhkt07JkErTg
xEIFes58oRDbwAtAPhKF6WqzKwZsjD7ppmpRzmrazfCXNi0ocjLOXVviDe4NBZbVhjOzCQyxBdkd
xbi6iyd0EVBaUxXpdvzrCypV1K7Iz2ZRVVXtlEjeHruxjR9YJL1APdlkp+yo164o3FAWDsFYMV4B
m2gcvu3neR4k5Chb7euLMDR8+L2edswAJogsFvZD9kIG/IHqz+hm8W7Yd+0YlcMcY9n1KIcXz4A1
uGMWkzL6lpDRl0X3dIkpffGrvuh8sT7CsV1fA/IB/BQjca71QzOdY+3LoE8GYkjsdJOTH6MTj5H+
4kJ/1FpFlx7hvcIoPwOK0s97JHpFavDT/1MKxaZ+qtzdCp5zvW+FlKJdKjN7ZTuI+f9NkgwyP0fw
VvzVNgluHT6rj1HpwU1x+1bMfcbr+P+eTa6MtcXd7Xx3pMcZ3BoBqUWU7j3/yrK4Ke05MvFxXnzq
9uJyvj+aM2rdVJG2SD77tE5rdrz9eQnU6VoFJonShFJvYsncvxueE+18C3iHX7Vjuc3sJSSaUfob
kA4YKg1QukVlHmhCE8iahohsBImPtsMiCT/Lvi4u1a43eOW1KuhEoQ1iHjeVEKvaW93y3FJHilS4
FMbOqO35jAK22iKwwmnZ/yEA0TT71G8P1NpX61RWdpDalb5TI81HKX3hilk97GqZJXUpe9pQyBeK
q8qsy3jGhH54W0X7SEmmJJWcJ+dDNhcJmWgTua1mZnRH4RPV2REZ2xb8HzuupztzdgWn6G7X8D9F
IVEBP3a3il7OJDem+bPmfpipl3eLBWygqTJBVZ74dlOzByouUMVOAskUisQouyszwUhWRbb4uiGi
FNXiibzIGwVYJhHGXqEaDHFt+JjwuyFZSrhGB/q50L1s8bZGw+5McqHrX6xoRhB/Qyd2sUoKWKuB
tQHURNMhn7ByNMsfKP0n/9N9/l+m1vVjG2Z62o4VkpvGb5YD5S26yA+A/wM+mnZ5k9NojHbQ9XRb
ohEYb4nR2QwstIbHOtcKowQ2VNEXUq76BQ5bYIa+muclvER1tpll5+71hv06biZ+7nVBSApNf7bg
4aHy9o6TMsf5YvtYMvbl6GvAEExTQ50Upw86FCvu3kPAnOyafDgBfhvauoQRNb7wX5vuXHiHcLBu
SHEnzy9uqYZzB6bp4y3vx/p3Gw9YxxnbLhuWJJfJF1Ls5Fqxp0uZ0x/XMGGYjuwYbVwullDI8oJt
Qp2IXDKJIt2I2AA0eoByEJ81jkwK9du7fO+/KzyMqUmOHevUXlPcDmX39xgKYO3iyMLs/VjS5jXQ
Fk2R1CfECQyEwTyqfYtvcr8bqmxy532/1m96F6XSeMLyiYtRVMzUeBoSPgcWhDGybiyT5LtmqJ8Y
IMaYXaPyN16qQK+CbWMSDr0er/939Wx/+EFhhRtOj8yXaj48s22oKLvEbb3jAlglYaTTkngyWZ0R
0C76rjEnIb5Qf3r+KwFQstMrpQkMPaGtGj8B/0Zc16tNyzG6dtOBP20UrUgpPXV+xhsLJpLRNOVJ
xzJiXBfcv5yOKyauYTO3r6WbhM07cjSlAPJWQB57mXYEVIQ3Qvw88V8eDKD1xyCUlIZ5u55QKNSq
vdKuUWxWb72CZCoRtcpz03vj1aq0Nq+MtkArX+Opk93DCm7l9mEejjs6k5aMT4dGoseRwV69Hvp+
1n7UlfFfYzzn+ikikMOVKsNqRHBFapXjY9ISvsHDnGtlJAHdoy4f2Wta/W4QRrRWidL9v5oN4bP7
D17LkYgwBI+jL2Vqao1/mHOKQM+/0j2X3gkAZ61OA7CIvB/WUC6d6zqIqukq+hPzlsVteKbUkK6p
flkKj2tTU7Y/C/SNlOwaXTTmuFypezxLh1fmHYOtsjeEpNYUR4qZKatlQqOXPNsPW399AZu4th1Y
srmrSrno/bjuQl2stL69i4PejxwlzPN/5pg6qrzg+N5fzm23brouLenVl01Jzg0U7bj0iU8pxdQ3
7ry8sr1NVk9p2lDxKl7sRUj1OpBsslfJUrpj+UFHsYzxzmNpwo3Zsx6rUj7fznSf+R6BWdn10+VC
GabmFbzKtgF1y8h59/Osghdi41TCUhtOktm8ViTZmpeScCbAo/jMmtGxMXXk97XwFqXb87glJK3M
fnDFs+UkniZj0Am6lXN0LZtvtNnkW4kbMf0c65hWSJsgnRxjJYzzHXDRvVq1YXfo2dMbbDlFhyT/
hlZAFy2UJLOA0EVDpcIQ3DpIl1SuoUyQLEX8u58wRUKhlWSbkBKKNDdX6mco3XPxnZvVAUvdf6Dt
2ZRaOkcC+k1i9bHuXcn40OdvTXuq/k5eOdcqYKpdie/2KoUgGIQjteTrBrSfGj/+44P83s2dtaS2
664bRuNigMB8BRGzsD2UK26vfHSsiyZba2BY5z6iV5Hz/4Drs0y2YuAHwMBoEBP57I0VwtI6Q+N5
VKV58bh00bJ16xDtVNbDakkNDZm0UeRVj0Av27P9nIoOZM9or76R3uBFukpVfJJ+Si5T20oQn+MX
uLOj8HWklw3MwEJKOQuYjxiikcHd9AdALGBjKE2TEW9HBnmANmjZvluPY9r6WTucGL3cocikHIKy
d5vb+2ueSV0r4zbehcLcNT+oyJOkdjQ8IMjPjoTjg33q8vlwCEVTispXUld9NFFwtbHjhmNMsyb+
L3fzH3qymaJqqWKhEDZHLFv4bE7K7vAE7EodcuGa/lJae3XPQpD2E9LiKU6diZkc9xdytAHESRkf
/IwLNUBuhpVPiZKX5QeyIn50bPTeAVL9bVKHuOR8ZhJX3S8IFdbIrWGnc7Wmw7wtE5yvu9LXIoHC
bJyjZGGirAH7X9e5mLLqrZf1voOqd9HwvR6dMZkmj217M8aF2bysAfT5ID4DCt5cT6jQ0UwWFULv
FfCKy0ouLrYTdR5cpDwtCDyToJOI79cQiALdQi1sdUzmHN3R7R0zlIhMIE/8GWzI5PCS5/+ew+DF
y/qEbxQ1KSMK8xGdpEOLjsf2kMTF7ZnPNGkBfM8GXKZayJvuB8DppKR2JNNhvbeeLEpOIehLYXUP
l0O6h3vXBBJqPAqt+v+YAYcaOhH6fCXMjzInZAogc/S/Dj6yDMC0CmJl0NJ31gDqVkn048xGJ0qx
unKma4kZ5mIxJx6mTl87nZvkS2BtvkVYajMBfTV7STs5xyuKLWMyqpWZbEihbPn99I42e5jBQyQx
tO9NGw8TgNyiHpfE/b+aJOA5HoWml6e8D49JyUEjb8tiuZzv5HU6ouy1qubVZuoGs1B1VEU9CRnq
w8pnRlXy7e2A2K+T0yZCnK+lFcRDdPE2lsJjy+QLLkdkdAwXYbv5ucM887O2BnjKigACD2F81Y5L
sNAsm14y0n4YVZ01KfzLjuSgtHz3kUGqdBKNA5G6zzjPieeVnf6SehzErt/RJmxDveDK5KlpABxv
N5igTefFpCvWJ+ykn2jr/LJAyrUj0cD8VKjO0AgYASmjbgGubMhJUq8GM4fVmwAWaYZXl0Cntwbq
DjxAnreyfS1kP7FACETl5irHOvGkUSQRlR7WuyGf9Pkd6wGPZktw/DOyny8KgyREFRDvX1GN55WI
Db18MhIsRG2LlgdPcMOkGvZxWwXKN1Vv/OABM1LRebohBU/GKpHSaV482BcEXgrlsAK1fiKsMFRG
OqcgpeyXHHmMX0KEhLur1+QbyFc00XGUD6Yw3xKe3arHyyDDIlrJgbDJuL0RsWq0rn3Bjg+fDuXi
m97XYJuFDlmSchH6RU88ihu6HJKeEWvKyrpsKOvuNL5cQMf0f4LiJfK/mkUTfm1gmFid6eZ0qnf4
Wyi7qdt3EYDBADuLqfrM0TIGNt9sjrtpHfbErSUlj4rCjRc064hddsV0A9vqLatW3bpjqLz3lEjx
aP54ePn0VCphiWGpsevY3TnL4QVgqpTneGMCAnfWxu4d/IuKPgZQrxcsThQlxd0LBFpY9ffqePXX
Fekm0xZYVu9hX+mWgsRn75PjzwxKD9K9w/Y3EjapCa3aHIdRpY20JBb4DtwQ75BFemQMFy6Ac4QF
+m2AS0KegtQwHh3PaH9YyFFPNDexj7CpwiQLWr7902+90VSrqAXxAgQvR2z6NqOShVPfmVHL89Jp
U4qxXQpXYH/7jg7UQhA3AnXrGQ0VQc8GClIag2Rvh3KM86MpF8GfJsJuOaOKNJzPqFVO2vZV3sEb
GwrFkIF/77lF2lO9zn+uiJ0p+oTt9rQsG8KF6gJ7FZipyHbkz81FNXudbofkI4umgXUhssbqgis2
3X8rZQHEojjZbxEhZiuqWvnYpSlWsstDceIHggWkiYZMDSlQeuPnpb0UDNXdmShXfU/m4o4QSBzl
aiozu291CFF+Y77TTsfnaimB87rkA3v4Z5tfbkRVKwGBnr9m6Wuq6aqFkRSn/M768oY3tHlN7nnK
6qN9C4RZHD1W7Ii3GcSfWAE3NTcL+r+I3rcyvXtyGG8cy6DlXDoDJpHYclLKaCwcGffKJ4zzxoY5
AYaqG47mxx8soTb7vzL83J5uoAvOUOiVSABQXRGo8FdqqZ8C+3OmS0gxje9CN5W3PWeCdLq2c7uq
OKEwJXnuvP/2fN3BoOwgKS4tGG8XVyuAh3OxWv3qMwL9LowVDif6FPj4NA2a9E4qycClkbb2PfXX
x9Duu/TZh77SwE2StuUGRoS3wbQVUEKuX4wHaz7cPghq7Jw5QFTKYDd9NCh2LS2wAZEjLq9DdZjn
iIrf/7LNiEAsMyirrax7fg4QIRTssV4Cb0gzxcrArmdF1MSo6mHMlWg8BVpNc6162Ruxrg1fVM2X
DRZfErO3LSBOBnIXq37fJ3XukKPGm++QCyqPBFaRGSp//d+gMPG/WtuaVQ/wYtihzkY8d8r7iQtW
fsVKD0VL+ZZ3+I2iF7jLXC0D6tB7S0WrjhLej3jw0TqThApyqNclhGkvyLZ8i4ZxwvtPnqeb8xnI
K7tyrNQ9FpSB1YsuxQ47RqjnjKXyUwPimPA4I9CXK2W2vtpFe95Al2PAkWhjcLyBuo1q6MrXkXHG
sWYpW1DNi/rwBMz+8jw7jhqk7YThD1aeOafmkAzpe+QLbFO1bYG8ruGIsOZmKgoCVRV2XX3x607z
Twm6iEnirs/O1t6HxHezIdMHjL9Bt3Bx5BgsB94IWnqUJgsE1DtnPN1pAAe5Hq5eOrfnbScLo45x
iA01D1yxW1rSpLIDUZDdBhiJB8rJZt76o5n//i1D73KsBII1DGv0Uc7kpUCc/UwpnTCPOvdy6Rqh
qbHVeHmBMGYL0S/Q4sYykEhP6piJmjWgVS6D4c2hn5fh96ecXpawE8lnNeC8ktSAEjLY2Yg1/SZ6
Z2glxWhyEc2I8Y9KdBJaz/UftoseKFNX/mz9F6oYxWjk8aWUQu5TRIgxWKHdXY31avXjNBoXGyxY
sapTeqx2VgKNgaTTfmCVPu6QK200KatLJZqI5HRz6MWCrwHUNExnEqGs9MFsUDMX49nWVWIEaOR/
1FhpuW4HgwD8dJ/7zPBBFZa0cguwGmfMY9A9CzMOX479V5JZv3o9hLgY2fPiIzMFaoN9BdeJzPed
X9IVW6znrARJRHYp0MKnohoG9EWSYrlpoQ1yRU3s5ywglNi2scdQQYOcQZoyEmH4CzCfs5RVjs4F
1yMOTg48JFdYDlT/FHxHLD8LZS/L2vXAiEnXe/FUzMR2OAgDtGHUTLCu/Stx3fFWKQnuTNi1ADym
8QEFlMqpsqz7D+DeZ1jCAJjgj4XZjbT0vqam1T30ty0GHePFoiaOSJeQl/VHRiZi6gC6EJ82Ud21
d1oOSRKy8cc9dnZQacfYbjxNI/URQsR347Oc7Wj2GMjAsfXAdVFcAWZQ6VtdRR+/uEevxOEGJJZh
ALHW8CBW4L6uxAP2yh/IxfqDYNc+shukbnZkwzft2KQvoFEUud2cadRbSNMFW6rXx+FPOYhS+Ap1
xQGwh1chc6S77RZWjG7xNEXnbV8gyI6fTIyc5R3UncTdxtUSAmInHRmR86YZS0H6OYkKYJI/hNgK
cxFptyxXI+wfe221R81NZCE7PGq1/OFB+0vwQyIId4yvqpRTO7fa8JHQwxAWv3jafy5Ku6vuA1md
LrVC1qXfj1bifn31EIJxu5/L5UE5Q8gm6ciwvYz8/0/SI87gKMwf8t88/zm0Vxywq53+ve7Hafl3
BGnCagz3PgfzqEvwDO0OtOK6C/PXSZXtEA0gK3z5fAA6pcb+8Gygdit0Jo2ekdkwDlkpG8dnTWtK
fdG2mvr/hOA7ICupenOCWDFbkr1nv6fYyP5EUYZuh5EI1b2H4Tyd/wC8KfUSmdNOATvYQaPg09uS
Dc1Hy1GRm1W9UCRmFw+1Z4YGrkY0LRan75OOvks2iVZ8h7ZsPE2MIIz+p5UmXxi6bYaG3ZgWabfu
S64PmOjlu+txcTHqLZCkJluPitrdyAYiPF9FBZeDDvVfrb75Fn/jk2Xw/NprCMrt12UtYmSnDYYw
fmvFaXGVPsphpKxT3/t7/sXvzHv0vUiTbObwEIm9jn1NzGnT4QIXbFz4PNvCGVmGYp3pVB/AUknW
/pWQkdsQO7AxujDLG2vSOQktR8wYujtsxworOlWxoX9T55ycYB4Ly8/xLbOhDqTCBQyAUb3xy3TH
wdsdjrNZlLWOjJJdZb6vzNdCmOReh3Qcj3W0Ik/bYxAv84u9Dd6hbJDIIDQfQSO/lU3poz6ylCxk
B6nra/3hQiqzuXQ06S9c+QEGIKvwX/rsrW5zyi/lJPjBzJc7c1cPsikiLAalDm12nJiL8mjiJrov
gJCCf2pMFUCOhA4uvCw+UTHkIn9jcoQfAfhHOpjPaQubP6InB4AZWK6hgY+m+k0xHZZ26cfAcg0J
RIx9vrL/GWkWIKOf+4BSbzEKP32nrvfEW2nzT9KofR7mA232RmkfEbUDhnmJNDwEvl1yQGJFTOhP
63xUElwQhb6UGKilOJ+YAj4HVLb2RiGlilCFN86hgpDcsHq9OjErHN7cDSeQoOGAT7GGak0YX4Iq
REzh5Em0Apn+3TLvtIQnUNwVhxuI2PC7wbNAbV1GfOFDijtHQJP/oXsJDUGOoAFj0ce/PofX9/+U
Qqjda84JleBVTRjjMyK1PpQw2sVKjSCc8qN79nULwmc8hFGCU5IkP+pZPQobmVdE71WCPeS5drVO
1CuXGFpJtts7ShTLOx4Y3EBi6UDqbqz4Y45lsCTK9zaGfnD+EhjcsGxRfQkZNeQfkORQG6NuDGLX
8Xns8z3A5eHR6w/oLEruEBVMMadv1QUF2yG+ewV49pXjrkU/oBlM/rsj//zhWfeQxhm9R7Ur+Euj
UWkLlWhjc2V1RDZdnxrXUfQIKjfJuP9RGtxKbWRP0D67jVRb7X7uVh0ktdbI29AuLT1k3BgO6bXb
ImFlXSIMhj3sS1RqSg2y1z84/UZVuJKg/7kkM1FA8/7Rvho4SECoUBmyj2ofPme2ChQLK7+/aHpR
jQTQakFMbDhuoHVtwF3ujx72iDQzeA5jIlbR1G7eoz6cbGfS+BWUGnFnNTKpasOVSS8r04+NiZ0B
r0h1dZJF1w6ppa2dD30tUUhgdsplNcSqRnF2mCxt0QuPp4mtaqTtsQCL4OnQJqi6NFGc+Tqaceq2
0qEBREEJvekyFUyvg/Chk067TJ2yTPHr1kvrsIL4blzeR8XZfggoFhtIabSAv0Mv+B+nURwFWRes
P+tfwAdcbkAy5EnmyzQiITclSbjDhSh1JnO7DY50Ktc825YiUuSSJdGeSbtGXAZSI++NsVP4BWN0
+0uzkZlHVUClcYuVy5JrncUWaxKOW5mYonHoyAelREF0LBQAp4F//ODkr44oTZ7FcGUvpyJacUF+
eUbCrtrll1gtweM/0hoDZ5z23nb5S9Qec6Pz/OCAg6UExk3vQDEn4yQG9JbwxhUWwLzHvUFMw2Uv
MUFaiES5cstvvo+95Y+v+8zyKYT2RxtxrClvRGOsO9ZsN0pMosUD7uPjLRI8ovCOpPrbIE0Vls2H
bAxlfCNF6dHEYsCXTWGPGhOZkeDqxx+zgT+RiPss7NPoNWb0BVITYCyQXJR10y/eTM3+jZ4UI7Kr
mo+ZAEzHY2jsuTy6Y2yHYZpV8Qt5c++KTaZlJzcagPnybgaCcJC+tZ3fJ8QMo1Cnuhr16M8GhOgs
nV5Rw2tGJ6U9bOnDcSdeXHn8dv2lTw9IAzodt4XxO0VgU9zZzV9Xy72kTauZY40slp3/qDJk3es5
c2xGPmTfXzyu6wySELNXeM/P6OAloMB+t8YYEzv0Od4j3AUdP8ABXgtihcPdqWAqcWvyuqInhp1j
HNs0rBnIxcEso1rTnnmiH7xrn1gAWrlEOVoBBMV4NBR/6Jz3oe3nCeLM/6sXagT8glNTve4dQVl5
088mD5R11xnvUltHGmfM5Y67WYdAvQV/VPo5aPbhJWcwF1d66Gq35vj3ru+v4jY4/pZF62RR5Vzh
QsCSZ0Nm8wrt6AdXfCu82TV+8sNdFbmyxIY3HiNcg0GD/nZ2fbmfQ6jLog+RtNk/XZEsh7c93xyz
YwLCP0dFL0ZGy7pNIr1HYBudcrjYByYvKTW0172Qat71PIdhgC8jtuyTD0eGKTCpLRU9oOPM7U9s
QqRO8W2R/5EH82AH1Pac4Mbcx4l32c80vJ50fCYZqr4+mAgGYoqlzUm+tDToo58nalNYxXxFAzcF
XMAZ9FB7GFw6nvKntykpq2q9ry72Vfp9jVVSszw7hKppOMxx0i30h5+lxEiv37m/LQrrrxqag2VX
Un/YaHkgOw6V9VHqAffCYibJ7AHBi5ki/4DgR+SyYTfWs8K7Fl8qsvGe7eVZ4ypCIKmj31MVBuR0
kMT+3KMXc9jauOq4p41j+gMvGFzuJ6b7HJ//WV1ZkzWkkfrHmbGqZy6f2F3+TlbTA/9IaX5PyRJG
rfyaXHmCZWgWx2Wz7hGcRM30Hzd/5g3kn8OgM74gXKcYFYVHTXWiuhBlHL3ezx8K3umnHpihBojY
tSNIKPsEzbaSL73ErTSMCm5r4ow7Mlrw/c2tG+NV9zOVQRG2gF1gzaGxrmlPoGWb+7/Zzb6T+ixs
CBT6yZDNyDm4y2+VGwp75C2xWo1B/EI48lVGal+FbF3gr2qWwt/jJX8axXDdlQEkPelPzuVkcNgL
e0IQJE81FTkChkCMOvHei7mdJMR9bYIONAepkikoESK+IUOOwDtvM55SDcWDvHcxcQI4qJ8u3ykw
mWqplTLCiOLnFBV3ris25hF4KNVs0jP4EZFtY4DJgHD+yHHjEUDxwh6/kiw9/yog6XkG/ECFN9vw
ZcSwn1t2GxU0O3zWjrnrHleqmefqzRNcwKqRi2SeRX5pWasNEhiNu/Hm8ixKjiqtEoTgQKtE/qfq
IGZSKNesquTKdsdmuTgt1Oimc11RfaY5PRB2ShMX5r4VyweK9Zgl8EuAbmDSN6gXvBKigRPp3Y51
Gus5nPJvCC2U2k9zhmlv5HZpBfUhhemQPjkaBxKFbYo6GNewq/SM+UMd8P7W0YTQJmKmeFZHTonD
+0xo1u+LuxkfiVuPGVSsNH0xzNfjTE8+97QVUCu7DwW2h9aOa27LPfp/HyqK85DHupubBXSqJ68Z
7XQPW5aqBAlJXmYPTc+XFFcbGWremMCmsG787QwsngzInLdXznm/jRvhrwK1gRoaa7/cKU//juRC
hcrw5zZpSOl3iED/EDSP4BMv6ePcSy4P72mpGQqgAkD/mPNeXbqhpScW5ZOOsH9hzESVPt65+itK
GFCGu4G8bRH0E4b2CfJ5HwIQc3AixHFeHUhOKJS59zo1QUp+LTxBgRV6nq3fTQDKfvGpxxUurszz
jeaCN+VVkJxDcoyDTi6Nh4wyHxVhCYjQez3FrLyaSnaH/Th78HN4y4I1BurW44K/MMKcLYiP7x+k
+eQBAVRHLxSH4w2bx8gewagD6DyZKeGM2RcDgOzI4Emy20s8m+3u+S+bLCCQeBo7cF96HNojeWcf
Sz8Uc4cScNizLgNr4+zSwsu/NQoW1fnMIcbAGiz9I6k+zU8ymBupIUsM0WjF6EJDYuoDyP/7DqPD
S4G10+3g2JYfe+Wv+B/afoFoojyy0cEATnJe/w6v04wj+uMx5VkCXJsN62bhCCCmmckg30+f1izj
+HFnz/MUYy6m9PWDVx/qV3CJpMHVHI8oHD7FsGP8a19O+lzebnVq54maIRJfG18IO91IbfFElZnn
MG3qYW/Kw5nE2mdDcD/iEPlBLKqIllHBIc/AFwPv3Vcb8W5EHNeQ+ExcacWEBCT8JZuO3njOs918
PiQP22c3iDhp+DqL3PG+XOLPoW1dEg7kOhd7wn8moePVh+PwW6RrypfV3l0Qj2rODKfb5TCMJHcg
SrF4oAI2yXKhildaHSCoXfGRCb7vbY+uGg43DEOmS316XlytDmsT8ipRCOgon21Fp/wUTGUfxyny
uI0+mOGHuh/mUPJBOnQDCnjK5D/0I8wbx68XxNfcA689wh3FrLKpjLnyoKuCMsWAsfIxU4uuTOR+
iMWku6UEljGEzjF3qxwyiVI5SynzkvoJXGXOPloB2NThHvEra1i6JQnzh7Fmkq6U2Cd5pWsv/u3z
72bJf0AOAVDJsTaRH42+cEgVmFw9pXCEproUmWLtEIvDuuj3wHZlbZQRJoDyEjJHAXzuov50FRd3
LzHWLTtIU4zCJBBccvDcxxVBOkGhx2COS0Ptkxh5rxpIcPdHkdJh6Spt41XwjKQ//6nUcXWvJbEW
wveDKWSIdovcUCGd34UE0Ir4FESs6cBNvCSztoifzeNaNS7gQP/ZLja4qAJVkXEdmFA5RvAonfn4
MHQe700HLbO1ZFh9s+MDaV1tKNoVFJPI75XEXjQmaSldt7mgl16lSyarl+SPa5Ph7qRHRdFLZ+df
v6iDVsccHdL3PyjiGSrBbsRxXEHpLXE9A9d6Ay5Hq91UOAWIShpWKBnY7n2gu2JkyRJfqa0GcUVy
5KPO65veh3nGnTXfYMczw5UnJtmYzR+jiC2mF15SQG3EqcQM8pi37K4YOkgzEDOqeWB27vkEYRpg
aRDaW0UvhcCMbQFtwCf+7zDiLJfo2sbqN+5GLw/mIBBXA9IWeHDYxA6QS/XH6QteDoYdtVGmt9Oe
lx6FN/c++bbGr6gLyKedHJMmAEffMd3fnSBQUTUm4JfZbfeun65oEEegESramkESu+0MzyBQsjLS
QDNXXxIWxGQfv2GMzvXCiDOVT6HwwJ/GwwoHmxhwDBWS0Z9yYOwa47quh4T7Poq3FiSPykm7hU34
BCypUZUX49m+s5vnkUxMuFwt/X9zzQUl2XgEerSR9WV6qGvYFyyyvpUcZiyd9Oct/OwGff4yP+ln
1iORvXOsebGNLPDSIQsEzGNfriX22eFgM0B2a9JHCt368pPU13OEpgUy2hBYhspHMEaHauklo/2v
pKLUG4ebQH5J7a8JhPYWyPRC5qYcngiSYX7lZH2oBijtmcc58InDIprEKT2SsCXHPKjehPUUz/nk
6HPbjkVfQJxfqF/N9yAaO/6k5DUY0vnjnoG0T+RekHiWf/BRCazVTZVpq/eGKdPtWckOcBNUQUbG
qtYDe6vu6bVMwmcs0qK/gDUWv2YB/YcqMqQ2DKXVx/YOokc/dNb4+z/XmAMJ/alSfnW3Ysva0tS/
AV8xwLo/zNb1YKYGUTTQm6A+sQSo1ycFdrGPBKe4aecq+Xvu7S2h8sQYWsyrLYurhefGRijCYr42
X5w4gq6nqb70336lQ1zRA1o1Xesn3k/viIvzJj5s4TvJ8Yg/le0SOc0oM76WHXRW5ia6nArm1F3o
VFXlamAsabehl51Zr7MIiLorXG24VXX5DZr+GOcH6EaQUzLnPnq21KAqcBJkBRnnXBOq6LLxa68F
MDVI+SwdIslPID228JgoSfRbDMGf4IebHxOgVh51vIZZOLZ7ph3chcuDHLfREj6EA83xtsdv99vU
FL1Br8iK7VJtNR/dDFR9Jt55377OQZ0KmEWuDlxYwyPu6e5FDWja3KoFsqPPnG2rb1F8+T/BRRpS
k8RbmZH8wLn1VHoYJWCCcoJcHVTmNY6zD14uzQufjHo4UZGG2OL+4ledq9OhLXlbDbo+82AqNyCZ
7RTolEjsOjlFiiSobueGttubPWMUVugoLVvBXCLxjTc9rGGwx9N9TVMEuKEn6U1UIrytqFY/jtDk
8CcOzNpSM7H2MCwd50epNbZ+ZG38fk+YTU1lBuzfge91u5EuCA4a8RWOCGIJvMYNCjXISNMZzKZI
9D9fgw4beR2LBPIioRh2f8L2Y6E9QAtFI9rfs3rx0K4KPsXp2en0CZgZGhLMNXq8WqgUuk3tNGON
hjcnX2l2LGWV6eIE+CcryAwSjRBlIR2Zr6jj9MilVLowfcfbxdrnsZfU6pjAWUD9u5oVPiFBPhLn
5o8AHJ7FrrYetDT5Viq1WlLtBohLmb9HRZX/QsPU2tP9DYe46Xck9bQGkLEQjWIemsdnfW10iine
X3mMRRayLbHHSEzynaKcGqIKGyPZBFuaEdElPhqlOKruEkH9SRwUbiZuSru9Vb7WuWd0Z9mbWc6h
CgSg9NbS5I2tEeOOgG6QobnXkqIPrzTkl5KrLdmgzl9BQvw+EmtOnU0Mh+mpeZIMJSm5QIck2S8M
Lf+HiqmvgFX9A2+a4K6kCfha0SYo3NSjvnzOa+bJ7ozMperUkNWmauEkQ8w4ZHQD1zqXhR6pY3lL
GKyWqvgiUrofbbmRX8aQFlJM4Okzdpa9PwqYe4BKhQiviVbRf17wKHRmJfFRC2qimdeT+8AaW9V2
KCnKuhljVvw+N5Q8JFB6DwI1NNQhi3y+Edorm41pWBEMkEFO8kvFa2/61iiiS8jt3IRD9I68vB6K
ME+IR6puTqen6UuMTI22uM7yHxck+HjxPEonBT8coY/TmQvhplR8xHgqW0SpwOZSq0W2DDSqkTNa
Ll7w/NJDIvx8ON/86fb8/Xxnl9tfBLPUc6clbfAneKeuh1f/k7VVlsQfhsBWoWrqQ7L4+gn+WJ6F
kFfVgiwadtycpkYZxwh/KKYC2bwgDeOgxfpfmLMxgDckbojfiO+s1DqWk1+ZW0hr7HMetNYoGlsz
cQ0jrVySfnR50+eyQZG1NwnqHW/dNfLgCpxHh+2Ftz/NtJRl2XOZAhSHF9U0u6GY5K3CJzg2RjBR
eV6RqyR+HyshqCYHNcnVUXt4pHKUWlEARmTgfPgf+lw8zTu0lYD+IkVutNVEfeYkEw+1xnu1p0jE
EUEAaIKQ6qFibDjCDT5dtk/CTvGF0o0IYstUSa0RfIF4LbOc1ysKR2gVFwpdy+NIgwN33jyk5f8t
dctybHiCRoI4KaCLtwpXMAaCXkOGiXOVdMXyf3glJngINujpMTubzMBgqoAk14QToyl/SQsY82mp
kDGPyChVLx6TYI0p1io5wjzbof9P+7H9pTQqQYSPOVk8Hh8WP0uWsXNobUlJ5aXoPO74dVXeuZcR
ukUaRfJH4W3oDQ6CAFkg3mwyYIB0j0RjoCgSV82AB3q92rmltfgUXg8nuOjL51PIAiHy6HyrAsBU
1mNyKFH37/9Nplnl/OEdLaCwwcJLZyU6QnO/fBKWI27buULzDcxVgGO/ijBCdnjVJIHe9m5+vEwg
BcsAMKNd1XrMt2Dk6EG/OHxxEQeXPuuTfDYG2Ps77aCvkrWALxgvDZZufZN77broUQ3HV9GpsXc9
PxGjukr5oE6jMJbOboOPJg+PbgHk0mZvAoEFPZ67XlfHgnZ6yAQL/ql3Q5Ep4cbtYbX4H7d+uGwF
NJCCnTEXErHB76ER/tYoqjYUe9swLfIs2cf8kJrJMUQVNT6u+reyiVfDbdKND2Hu4BpylBGUGzKJ
jDTtvhOGouw1YQTAfRE8CVGE1VnxcyoCwMgrpmZPZuk0GOkKAGVIoIxl2H29b9LOLFTjyJgJKVWR
L6Xhho2O7N+21k6DGD0R2P7kSE3+pRbRBWZM/s07JVuYq+A79j2beCtGTzJBLRwHXENTpLOo3QO8
86T0pih9IMvSVrNjhwuDJXRxjoP4ihNJRizVTsxstd19yELX76dfH4+MygWnijU1KwjRUNIgEABk
CwXPHVFd5EzRDa5rzw1zSkpALsiD4e1jzkLeVAv1uody6GHhLEMR7lUkmHQFksAzok8AoPic0BHm
QzP1WNmxophcesZitU0tkhk5Yalf0a4SKoitoLrLaBDQ1gpXufHOkTRB5BYtMyvaK5AETcc+YfMl
A3+mXqaJpo7N4bAnViqRtjQC0Ggonel0nrxhlv5U/5bFFmDEMH1zPLVccvrO6lq8n5bjbUWrncIJ
OSq/JzQ5GnfnE6iBxpam86i90rM8jDyXvLMTKBaFcR1y0zkpnt72lQ2lz1le8Xcmxz5CGfX8zSl6
YF8+dBtp/uItlzaubMejTMF7M/hmbJxoKcQJivWDJT837oxk3vRoCtaIw8qdKvY8EYq+FAETwbiT
pLOoHxQO39jry16EqXZtXLKJVBVL2jBSPUj6oJRippDehKKWvBuebg4IM1chFeKmheegCHJDZnm0
4UMYzBCNEPldJpoa9xUBK7FtehulpN0QYC16og7sG0BpzHRn2G+WmgcxEfBHv+/SquIzf8nBgYhP
Uo6lK3/qPX8HeqAyneZ7kTAtmPCWIqnHBC12Ijx5XNMOY7WYrRZWGF+f2Rievp8pZwhlokTaj9CM
GDRcwjTNkpsG732m4VD0TPxmYyZczO8CizLITi8jRipSFVl8w98rilSxGFuSRrigWx0RHpUEvQKP
fttHEy6MzkK4+T5aFxPYtM7vrMRy1A4tpIZUQzJJAfSzjR8Gx1/AAhXh/8wOZ7wkMwCFhzq4Ou3E
oCpJqflb92e4zx3HaJxoXmL/4qxFuc1AxjJC56lRVXwlwA3h5BmuQC5yGDISy15MgCtwlbCBNFUq
3s7myJZqXkf34V9iUweZrtO7cTlytfIda/i5vdLJJHvfRGpVZq2bNkV9gF3s+6vGWG5Typ6mXSQI
cKMTbwaN1AK41MtLdlzJlBkNY94Lel680wbLNJMpciaHwwZo9zdINw1EG8VUcT+9ZI+p07AyrQj4
PROhC7pJTPz/5mV1rg7waCCPhkW3SgPPgNN4BwvaWwMCQYcrXVGhjp6rBvZkiW/vZMuUmkE2noqA
LDTM/XNJ0sDHzJ4Wjq2ieUzpZUTbnvQNIn6l16kRukXG2908bkEW3sk4JzQ/GU+NpYysDRFFRHhf
+cl2Qn6vb393kQRf3RPZYFxEb8a5zlJaT9lOq92jpviIHZmdpFKE+b6XhHdJK7AkMgX2eO1paN/K
ab+TY0Me+v6wbL+F2aSQUWUVmPELlUP5nCsdRp2U1FTe1gONTJiE9bx4uOOjvqZd7nApHoraMBWC
UqbekVLlpQ2wMlrqSDDMNYZ2IANqRR2xs/1dI8vZmIOnn42kvAN2BmKcPwP0ysCs50FN0k8Ycahh
N52jn94oFX2mVkyNw7I7LT0jMPTlowK+qg2Hk0I4I0ipwQDZgxwLtjn0uc2Uv9ey7sqxnoxUOmOR
eAY+OC17mkEjfeDKTLXD3Kp/YqoFym61C0Vg0bvhZX4MZna1qKfmct2w7rieuBg6VsMWPGI5dEXa
zZ805UbmKD957KCMenzUFymjPi3j9mDsBv369FnEMVx+ILL9VlIDkQJQmKEFO99rAfBToN88uQRf
DuLJ9hnX3Z9CcVePrDmHSC6eVtpI+ftxGfvW9vLKOmmTxK4WChWeP/psMB5wBU0pQiMK2r0OB0pI
v5wiQ5ORYXuM0ogZElhV3rbFm7vzwCIDVvS1f5fJlz+SYRxT/1817GNIdUC/TFwK74Zlt0l0VDDL
U/tLXQnCYIRCTFtyZhlcqx7aTjoNRdSDaFFhNYa4RBwaNwflVZVzn1jAzRny5+A/euKxcdxale7J
fsgDfluSe4SJeljk9ppovidR94k20Ns22q6P/yLNV7LreJxQAqj40ShEUKJFhS/BEi8rzuefFgUL
9hr1iqh22zd6jtxA2xIsxBASR3TfHZ7zC4IzMsYUNmP8PkyBaQNqvBzfc6ASeIv4J1F3LwG3iyt6
6u4d6aG1DQzpCs9W8kpdMLMzO+Fo1sYkU7kaYLfj30q3Q1t8cm/yI2EdRxzwJIq5csBCE2cMmjup
Jyd90J+7KneuRg9cDo3ty25IYRbWIWY/5eAcxWMnrJ/10xW/UH6gd+V8UZ6LjnQNvQLv4bRLCnMQ
MEYtqnU+fs0v2rIplIhAQ/6NYKDSo610L24jte0T+OJ1Xhu6lmkj5Y8EJf2i/T9RO933r4kYfFs9
s6ZP+5unotKlOYqby8s5TlIxlGX7UgmgZ1lL9d+zempJBOcbC2JfIzCqshbMhDogu0tkKGNl6cIX
iMHY05lb4kbcGfjIL75n6FFAt9aJ4c89a4dUjjmqDX+wMGE4RBwXEfN2zxyxvQ+MrbWlUdGYqz9x
Ci43iIWs2+iqDJoV68rW1NKmYdP+53Us+f3ry9r1I3ca8JN/J2/FJ6A/1KMRwU8xgwoL1Yy5j9Wu
FvWvLkPH7E9+Kpkv64q6282k3drR9djHcJqmQCrKC8XXZ01g/1k1xtC2jNQ91DpP3HyfSoZzVKyd
zI6fVxaf2WV8s3Q4IVlAe257yjoKgMVv03ICwm95JPDPFpzA9jGpbMRTCTrU0MTxraxyFsk7qKWU
hIa8XrItgyG5xc2ife9d7vTXzkZv79ayPP4nNBkGsdSzq1Mltimu21Ur4/M2H2/PtE5SJ4pJkrxZ
f+1P/9lJx3TwFFJ36HtuA4CDYNCY05WKOMhXQWVP2YaGav03pwpjQzgadLUP/CGNQTHBItSO/s56
WhwdrH/wbyBaOYD4vnH/RhjZ0CyPum4HiF9oipPRTNFKUPbLYW+QwOjJaWJRyuSN+Y1UawbxeuJ2
e7ETuXwM1b8OkLAz14Aj4QTuX/vaoLVa1qjBRIPAV2InQ1mEN8dksNkJMDsKQJ9svz4vqIyfn5RI
kXkgO0NtKJ4vQURUMDZ5jEg+g1u1wccYT0mrsfTWUUAXOQdly43Ef+Jpx9SMOzNvQuZkmXH1SGwK
TqJ0a5lOjWiMHi0y2CtWvWKlu0fbZRpZhbNucDBQn+3OjDTcJSJP4qsJ3mtGMD99OsSxWvENTKth
Pewjqx6/nuh/M6USqyUDRtKx63h6t8JArVTEYGeVNlIhKuePrFBYRCmwd6cO+sXhTdgeQi2zYiRQ
x6dvmtR1kfXwyC7NS+aeKq1nfGijYy987bl6fb0PXkfF6bUOSf7SuYfr+3sWuKLw4W2BJ4pMJTLb
3WaiKKxxdMexfOPPl/zbSZMv9gcPGSQ3tLOSAeVKn93bhCYQCIIuSjPrTpF20s0BbiVYXD9XRdPn
zJ4HfeMX6EMTkL8CMow6Ld63pYB2vxTI27yM8cJHEW9jxdqOK9Bb//GAt5kRjbLtztmC8p8TOQ+u
OV1YLK3YUHqYw+5yEFmjnKpUw6T/sv1SGLEmW0/wyF4VGjbngcU6GbRfBDUNQI0QKJuZXbPJ/3xY
p7wZvZardgyx7rMl2xQlyZPRdn3VfoSEjOo9GMIbM4zlJzpDkDLd9eCQpunFEnUwmgFYPob0zfXB
lSQSUX1N138TgTSo00ebgbV5UDUVRT8eipDz73vGi8c3Lce6PIHG8NumvXDHIqPPnvEzBtKv8+T7
/RiBA3FM+Uagp6bBaLtmHgbI2MmiCvfoQ+U27qEPEsM+5xTT9IKcyWfke9aoYAhA2s24Mrp+QKm5
grGviz5XOHf7iZ0wooxNtrZKjXH+sm9Sfb3zoLcLe8lCoCdNDZY+sKeyE3DFlvea3LnclZGuZNDk
joGB8PKq9WE1jXxbgvx7ZxwG2nulGBBwS/gnaoWpz5QpXl/r0iK5NdDmzg0HDTL9FdyUNA8m5Vb9
/Ffae7nJOXydvdQYByDoxTIm0ZzBz16Q4UFSQ1CNkNHliyaucgjC5byk7DRqlck1OxgXllBNvDOE
LQsz+A9u+Lt0RB+e7LLxC7kTwhZo5G8tm/bJiIPjcSDNZaCLgs7WqC/yeLVvLoyn46W2y7/ykLPZ
m4PATDM/rrS4nK7F+g0pv5Isq4P1dY04pIpK2B5HmZptnYHux7996QY22SsPsxo4vgxGTcoDG8Lc
WiEkIbpW7QFXk92fVOHahGjeXdFv8CqkJjgoroQDD7p5GOWyVBa/hdZNcFA7MlhVxkC0qoKRegdz
vAqHT2+MbcLHOdWjDH53Fzh6uCv2X7v8wRSgNa+boC+YmzQPvXcx/+zP/1itDjGLqYKTB9M/a3T7
Zr1AXtL6cAx1Pyh+TTKld4haz00Rm0a6+uikE679fIzKFLCY8Baz9LjsHIvX7Z/6TD3wrnpgwzxf
BW+IZRTnJlP2tuk3Cq6C7Xo6sFKLGrkGEiHmBrtCdl2WoQ0p9ufdH+tncw9gY/+0dWw7gKZsgL+w
IW1XI6R+KApAA4S6CmjvbpZIkM9If4P0u8Djuqmc09gD91hkViXFOsPiCoNt/GPgoqGLGlSmtnPL
6BpnJKjAPAMclJ/aMam9mC4/+yPUu3efjajGae96SoRLDC08OQwVQZcYa6Oauu+9f5iElvi5EH2I
DbMNZpYT+/BfbvLddbyBcSCkgqAJVfQX8nAWoXGgknLtLKX2iW+8gOMSCiC5gXNk5sTF9/bW8fBA
GW3dmvURy/FIR/LEbXK4mxsfBcH0R4MfM7sEol5eG1dFAJZBpuEqyYDRlTWlEsN7dsPymA/9rzd8
IDDv8eErf9otQlwJ18p5vz7UVWwm0o3VU/eU8zkmR6DLsQJ4eGvtq8lxTF70KTOwIT2pzjSRyBGB
qlHOawtaqiqp4zGDYQ76IojIq5ptFOKN8xF0S6JUaKExGFuDc29aXoJkzU72LGFOl5NHSlsyNuYy
9CbEoBnJwo7cRsCvbx9CZs3YDI0nhd2a75/JhfCt7b0WzeHfskfMpwPJXGOrcfrZW8C/xaGaQH4f
iAM+pwgu5BVMvI/K3FZzGGjIy00yYsuIrewP552QTNNp2j/fH8VCzet4GU5in/IPzT6DrAToRNLl
mQM8IgU+4KS08NtLfjBsu0KW0dmxcJx7A/DVU9wq6fBlwmfLtCXAcSyypd6VzM1oMkOnSbjLE+mB
cgru77rhMSJUmI2ATZhvaE8IQbIvHMyqz6XziHU4TlbZqEf2DHyU0Q5yVZcWJs+3EjpsanNOHWBH
HuLwRXuSKM9jadOBEl7H2Pc9L9qYKj0YeuZXXtoXc/yLAjt+IIOLE2j0H59ZBUuwQMDsKy4ZisiF
Wp1rCXp4OGkGZYeAdh9YFnrsv178ekgBravk5CHviU8t+grPi5Zd8V/u9TVFpKniZrnX1c/NuNJF
TCraQKXZq6jnpFq+7aTInI00FCY+cIDFVXczr/l+UClwCr/GLHYyyuEBOR4LjEL5awltTtA0w30i
WZo9yKZ1+1qGYxh28U6TiWn4uWyH1+LXAYls2qo8JxwpbFbHKbMutt2Kf4iNqniDSYl9kTX4lS7P
G2PerEObj9mM6Q8hi+xeh/cmI6Yt+OIBYoiAI0zwWLkv8riuYjtpkJZwXxKExf/vO/RuPvuXk/p0
Z5sMPuqhT68J7gsm2Q75kS2E8UOaGBRCkayfovW9JERt+K3yjpiuqs04OIz5+nk8DZOclLDbG6Yu
jdnLIXZdQuZ0b/eSw17F70apcplQ3FkgzkzfGESvBQtv2g/S6H9myQ7wOGT854xfYBMImo9xLUNr
g9b4J9K3aqV9enHDVCTOsbBj0TPAk5Sfu03u19oUTibUaSxFhgsv7QROx8kwrsyCTtaNZvo3wKY5
3YdoWeAtXMPEFrbvTyQr0GM+8K9nOQ2JSsAUCV5NYIAHhHXJrKjodALuKY+WbFGpSrKn09DfIwDe
JC0U/GVGPLuLQlziknDvBnI51xMxqCD7a2f3qHRsB8HI0ePH12JmT2I84lcOlvvJaOJcJe/yW627
FgHHIPrky0U4AcHpUKtqpLBCEiA685x71XM8bhkqFGq5dhNqpxooYXqK0chppMybaXyGeW0iZlKO
saLWDmmIhZDnN/Mnq7jSngFT0OvhqPxkQRua+FGjaSIGefkXXx9gJV5nYp4nfhoBTRbtwdDFpROo
MkIvPgQL+SrSdIXdfZpwYVjkQQI/eDQsKOMrjdpvY1YUFIFdwBzzMfYUQPAU+Uw7YV5qIhtWdLSP
0EKGnTFfdqK7wHnRe8n/b4klIGCaxJ9bxZ24PDWNcc/vj9wp5OS06PF0tp3ATIScCoKCBoyMPl2f
vgmyrIidofFbXDv9CWSaMFzPp8b+OHV/HAtIDNNFRQ13MxvOBIcbDAnkwU7xLLliPMCANnP52Znj
z3k0U0JiOh+0fXv6P59JPHgb9i6HwV/gQSrZSCiPTwRW8CgBGZytZDIUzLmni3+Wp7eSp5TQOfZx
Zez07F71J3eKfv/mB3reK8A5+JNZBVs7iMaaKMI8NM1GTROTb6TXQWMAS7sJmx7OZIVOi+HoFesI
/G/CbmW5lxzvF1YvBU2FlIbDf65ZhmwcymiO3DyDQLJ6JaSkambLZD5O6q6HNclnk4yKnHjdZ9bE
tAaTUfEqXcoRL4qCm0ZXnNKt/PjOWlDj68xjJgGWyI7Bc2vIReJJGoFPIuUJA6z6WXgWm0jvIGFM
XIcgS16eo2JzhjREqBnPs0RoK56Zomi10Mzxfj41j1gJT8Qy4nh8YZ5xniFGtywAvo1iWGDv0Cow
R5q1OZKPBnbUuq4X1eh523SXP2DGX1tb4GKRay9bSW3KAeV/j0AMmHwXmwcS90MUaUdQYBdL52Hm
q758JHHkfwxUkF98DJUFgag8L23k2fcpnvVVAdhu2fUZ4Z3cpnfRiEqnCHC1j5YBf+kvPwyFLRQj
3G378EC+2oD8pKhzX1dWOxAnp6b0zpEo597zp6f9y1qDD2MdGrz2/rJ/iZFoXO3fIasudpSFfWJI
yTcpwWdMjrRojZ/RrJhmUXBcDMfeBUwL3H8jqmlgJFEWBRWR2/XQBQkc1wZTZ2X9asFxLROXp0Av
p7Let9m9AMv0aPTINpPJPnNCHBm1jKT5paTa/MPlJeLWeXlyxCdy+e6RuQV9EnTvq+/BKi0Bl+uG
ZGty8sAglyMQ+UWeeWtKDbqtXHRO+smuBPcBB+JRaz0UvJLPTlplcE4fq+kBd3CiOe9bYwSwg3uv
1p3jZVG03E6vyFX4DN2/w/YIPE2e0GiGy51bZ7Ms0j+4n6dcGoG9n7BJUk9t3purorxTYbORWHdt
TucRo+2XDkrfw5jVScyak/EEm6E5PVW6LlDLSfopQB09GPzpi779rUZgnF7IeoChSiWKhs4URrgp
/uBLwBfOtDhS5SZVRaFqAZfPrTpz/pqHe5GvAU/bNngFEr7+hecUszKuoLv+5IQUk/FRGHWXMrBi
ZsfBgwBHhclpHFYMkG0CluLRaouLMiF9rK6PwyRs2V4JWDRNUFr/BJnRCnoR4Siz1u/hJC5S8BDH
zMfVKch7eCua0lejM2MUA2B5lVK33td8yub6VjyGTtP8KXejlCQJkTOvU8suMGYo3kFtP2HwK8OP
AiImnz7VHMJR5GzszimgsYnWEyqgWVzGvnktifkbXVQXceWm35MhOgVEmEFH9OIERyL63c9gJTyS
/n6nKUWIhTIIokXgqup48FFOOFjPhu4WDEECkp93NaOCdXl7Fr3/PkM7lccajrJx9wCyvfqgT1AZ
LLF4LEsHq7Arj92MBNMsDiuAnUWPqpPc+rziUoE4Ngl5PH0FudFiQQD1xWQMwyQOvtz7vRLgDwE9
Mpoi4QqNoKJ+yj9FegNTuF2zI+1EikUbd2Fs5jPNHDHs4FCssL/6Wblsb37T6XwTItvZmCfv5Y1D
bTyLObelazMgABs6T7gFLjNzr4Shfkpn/R+jMbpQYMCph4Em34qqjofLHodG4XFViP/7KkIzPE3P
WbCjqmDduotfnMIZkJ4qNUgcWEYoNZlOaoKECayGPJ4MDnfG/C50P84465PFecu9+yl7cl7V3EmB
ujE3nZ9wpb8aLNYaHCyEmbCqbXrFKoR7pU31Hb6jcsARlJgTNrbFeX0za/eAPSnSeymN9RhGw5CM
1CgMCM9qjdm0l7bLBQyi4QMEqr8v+6am/aGGFtFV/V4CXfcqAhPjYDFR8qBUZyFzPMaOszVRXJUD
uwH1aDB2mE98LHmiCmna/PzVrQi98I/Vii/vrNncJXc0vV1i1/o7ZLxIN2U3sqVDgYD1z5lqOhwq
yQ12HFe1aaxGPlkaLYq4dAYvvwLmiT1ER06lCOSuVn5/BdPOg+svjB0YlL1anoISLXXWHC+X/jCX
PrJOsgu6Gl6Y6TX9ekW1or5cjPySN2GFllgTD9fIA2nYX58ZFcOuuXDCB6/B34LtxlmxWJfphGMo
STjAI1SnwymuyeinrzIOM+LHwilCN/Pk2QY0BEAx3zQ9CYaQmWMjjWvaCQlVeqTImZKcpC2SCJcZ
Pv0Vo2zkvmTc1HaooqVnMaGvQztwK0C06hAZB9dYEcSAVcf8CVM7+2sSGciT9fdrOqfX79/mYXZX
U3WtQ9dfhanafMqz8QJBBVXbTHXX0igkpWWNGNjzSZMYG05kji5EkHRz0K7PwRcddYfKEYJvlt21
51Ouu1lSpZbfnUVAMsnm+Qp8ttVF/R2Gl6Tf9h1m/hN0h8ogPew27sPh0yl4EYybNyci4EDgoQHg
kawCD0MwJ3HkdzLd4isw4KEy9mcu0J2xQUUuhSqz8EeLdzYbBk/K6JWL8PaKtm8kPdZvR+T0FJJ0
g+CdPOXxBBcgYKF0Kd3EIOdmWM9QPmHvqeQjnLtY5nBnxdHAuel3q5fRDwmETdxyGbnwRO1Y4lHh
PWox0/kjZtBCCA1mfY00qBO1VFTChbN/C0cGOWh1NVjtqe9K+OTQrWUuhbaLQkLTvyehs5upiNUo
Gsfs3NB1527439tuxzM/KeXN1wUcocfxuCPBqVdL3J44DAu+tXpT4RsDeHXIXZrhgQtNn5vx+fd9
PfJcPEdNu90ru7wJmpsuKtt86WdCmhzg+GoUttJ7x5enYV3rSqWL6nDybauQSi8HaJVUWx4UIY/X
8yYOuKIwpBxQw+97E0d1JTi7kx5d2hz8jN2Jml7EvKWQzUI/y70scp1IQsH2XaLK2BmF13VQG3kS
CVSTm/+oNTdwLzeueRieuOmM4SctAorJNYFAMT/+OqPEcaLxJ32nbIyBj+3w3kPRnd681FrBoZfB
FcXq6P6QNr7ZUVU1IyPB38Hz3dAlmUe0E4LY/yhcLeppdiwjnEOinHyZH/1xAuzCdvMLOC/g4ViM
p5Vm01Bmhs9LJB0iG6W1u8owDOCh+gTz0TvCNHEz/cHcRgbNS7C2eBrer8ECrALV9HnDG0fCtOHI
MU5QZxaaJKPWwEZn+AYiPIJYVqDMK5ehEnIxQw6vcGT9/raNL1W1cQgT+K4PI/nn4uj/AnF5AXNA
yugFxmZM461p73hcUVvf6+oIrksDFi4JAbBMS8pNZRclXDbokBzcgrUDznabLguyiWMKDAYCwFdA
3F1uweYaFN2gDxtXkglIiz0VouBZJ6eucRN2srr+PBfxqDLF4YVUm+/7lRDS3tdSm2YQifepXO0k
KYHOnzyENRq8HzTLRXP06Xt+ok0YEpq5Ni9Ob2UydHqtmRB71onJ0z9Dg2vVKIL9BBtcEcVnbUcH
ncfdJb8DO7eL4Mykcz+CDwmouj7d1eCkBwuGRDKGCOnLK0TKlGZzseWpdmoqjhl9adU17gp7XoPB
Qzie0fbqcbGWpdWMxK9R/IdctV+pPv+7QsJo0FRfBPQuhmwJxr3KBDqMowFYocGmRMjCdnxbOUxL
U3dAZdJbHcpTJ/l7rSeJ0JOyWLsN48g4vALDAUdk7tgNguNZJ4e/cHh5iT18XszbNJZ2bn5OhI4B
cmkHxCaRj4spsOAgEgDrE4xl4MlWcBldCsLUqGxEMO/Jq7mLq4EWsTwehoCFYzXwTkQf2W44Srk1
9iFVfey8hR8yWl7cXRZQBOw81J1+S8fLPMIeMqnDpVtxGRvAB3aIilTp/MIsfwiBAurPtP92rVy8
LlmnNGywU9cpTKsjf4pXQu9iZQFLfPNwvsx+C+XTT3TG9vXPJSIebqnSUZhon1Rvx/cYb0A7xWYM
87ZcE/T0lTMwtLAVSqQKeKAY0Ib6nABAFFAfuyp/eii/FOHVq3JlwVIaAvSYf5pGf8ZRE5jWS74S
McW2ebFesOpm/UL7n3VyVc4TCFm82/bOuDk+YFl7MNlt08QAn51F67IXzjFbetu1zfgozJOp3jKL
fwX8Q3i/8G5kjpDZOkoS9qmCYFlt2Oqr3gdSvoxgsla6iBnWefudN1k8ZqRSRpO3GlgxOMUFtJpY
sBqoWCUUe4s3FhXd2UIC83LR0uSdVK7KmmXdOsGrZZcM+1BnwvIaSLQunJUCSlg+q9yydjQ4dzYS
zLmS7Sdzdj/Vvusuptie4IwrmCK7vqizEp9U/ANwx/dY/MsmBtQp8qrnljx17vQVnZSyshcJ2CDa
MncsdilRSnIWTYfZZ5lQ5rvng7SG3yJfTyBkFuYozSZoEhHCrn3SbbRQmTwB9oEpNlzuyyOI2EMA
PSuVaQjiiv/y6s7xRYPPhfotPmSrhQJQ/FW+7oTmF8Dr2SEB7No/UOObHFbMXJYQaGwq/ohrC8oB
dvW9U132wF5WT7FgPKs6JO9Jhbkfu1+ag5UuRKVZe0SyTprbH4vSAqV2+R4H1sdHsmiRWVggicu7
s6vb4+lcR3okdmP65krFUrt3R77jxgQnTkUzOMMwQm4tQFtKdDigomnRqd1XaFGhT9PVlKfLj9M3
lJthD5efdpl8CcqaBQc0lp0MLuh2HI5ch5CJTR13GPn7aEzqBIN8nB3gfvSUg4LqN0DvgPYFCTx+
9wzcTdjzuOWpWWUys8anewp1Q93ihJvHdkZ0qCgKMWya1ks0Z4YVY1sPDSMbYJGaB/TcR9sTujUB
R1g7BCC3x1zZuwA1tR3KFjTbv8ceLwfayPIv0h8fSCjBGiGTRbX0ZfCqdwJOmZjwkFdiZl4Uyd4K
5GFNNElM2L2Dbu0OQdCdCM7WKa7IZeBrtq2gLjtqP6F7B1Vrk+X2QZWjj+nMiGtja01hCDbXC0e+
npD5NGQ3SHNZVgLmorG1zO+LndGk2JEloqKX1C3NsKcHFxyNPSDJk5ICTCakjgF7zzzzWeQFIBKc
cqVNZgMVE6baAIzlTvaCuYcs6rv+qlHczF5+3C88Fc3qnuT0iRBXeNC8VDPynto/FUFVm+KOEB2d
Yq20ZsN3OEleOIuIt6yeC4u05hhZvnysClCpEqyJA5UtUbt2EIVT6xMn+V0eab8QUpU2u1yIhuTA
HhbZJZV10MR69A8N+FoqJNsSHMAb4sVAOtiMMPzisN2A23uq0+lRxZYtKwtcLl2S9o4PLbQPQR7/
+CgW0flJJezW6EVnyrtux+B9Cm0dMxs9KB9pW0U/NgtK9yE2DajgQn2UALo7NqGG84tDqCrg3jFb
WjwtGBRRYe2kuEwHW4dIi3C5rvKfGTtOUQeLWCW1mEx2SVPDbbJSjoLefGYxrYzPBpu1TkXzWdkk
RWA8ZZDIKcBtj7OQH69Tl2+KaK9s7gftQTBXegUOzICmDssBTrzXf7RgqZw8djJsjOEYNfGJWRbW
t57/b+f9YLupRU9spI7WXZ5aAukyqR45zIssycLHWqCB+Kneeeb5gVhBSr9hM8tz6ldN7uN+M3BV
BtEhbsBDYOcDl2XtI9Jlnea7pcutcbeSdXM3ZGkBSkOk/vY2FzoyOHGAPMPm9bgawgxT9elr3YgA
OOv09tg/IzPV+T+07PfJRP49oOYarEfNqRxBtg2wV+1iVjYjqf9K/c9Ld1aA+x6roDUslnBAO90g
HPiGaN9HH4yvRnn8ezMQTB6+VVmrXgmzqcuSomSUJjgrV5b7HZri1f/X7EomnGJwpAzNKHwymnaP
bO1lJntgK9lspR+1yeHqs0Inld5xFr7yhFVuWtRyCuTxJ+6IuhSqRMtzW5fM8PWR/FttUOLvXj23
hVHHZQCQqHai3h2CLIm9RvukM35yQnTqDDbeY/KEkRSiEVcQktzZj/Vcchfb+TCkN5gKN7SaMsjj
ly4Gc1l8S7UP+ZiwYW7Y7NB5SSvyjv3TbKNu3tneOD+WxaLuo7bgvG27IPgFJJo/J1dchETCM0w+
QPedX4s1XqBUYiTm2okI6JYKYYB8TOx9N7t1DSwB6H5qfcx92NgQNCJebaKT3iMzHCaFJVGZPzve
tM0sX4WJ/CnJ78uVAWillDzaiKZJvML9Gk6H2kiGtiVD5IxCoOwdCi0TSkfze0yCmgTwKR5CjhV3
6zkLO6MKvw8y51mVlZoHCHU5jOWpdvImJ5Lz2W0PLL6PG2dF0vYu0LcG2Ggyxkz1XZfjY3OB1Lt9
WVZQyjUi5ibpSXRjrsB9YQ3/GlmC16CI09RPufdvbnAGsODft8hYsGrc6HDuezTwZpQQKn5/BQKL
1D93EBru1QLF4GPXd4QMIzAYqBIN1+dRIbrlAD4Wb8nCo5pduacP3Ziv+cY/I3FFQSlXv+tZQada
pO79Due52z4d+dGI5drpnNmpyLVgDqe5jhDmCljUo+BU+NLM7ovxXS0l6wKZ7uSUmZ4gDyH22M+5
bXr7p6XvIOF231Do5fjHz6TzSdKdgxgRXcfbc1/SIPLFGmvR1qDTZwKT01lTr3ZuFIZ9OaOxXcCx
ejFJ1T78UI8ostuE8IMs1CyBKhYsRcjMwY/32xJkSmqj5KNs0WUUXBiFjyfkxglM2VKxe+p+DtaP
xzPoa077qCsasmnAOa1tbJ1v7sphMycRAVvNR5TOBGEfW80jVaPd11FsP0z9Jl7uW/8BFzB/YlO+
mg3nNaWduX8Z/tR/57C/bxbfykzOe+Vj6ZFxUpysldIdROW5zi/62OeTcy6n9wiYo92uPSVYjfhQ
apjsCLUlc4F12jANvGag9HTH4WcHOsofBiEhlybgcM5PX3IZTeQNwRnYqsguYGX7cgvC7OWI6zMZ
HvcIOd/QOtPp7ejJ/4LKlu3MqOa8Jvuf/8QNqiP5tkFxHLwke49IfRz7yRhFq9LS3O2tgWaUoyTX
InFntxoMbFEGZSWvj7lw7EKAtECHAtoKUMxklPcxdVs3oIBaRlijSwRO3LrtfR67VRMgrM3YJ1Vp
rLxl/29Amq4MN1IAz7gUkGL3WzZG047PhnLx+CNULz7xV4btQqWFtel61+DayWUU3Vq0uEsvs/XG
57AIWJ2uUAyaxz76CYFvQct5grkt+3e5w2ji1PI7H1k+iacjEEWupDclpZ9OpXRihkpQBJKrE0Bv
IKNlYa1ep2OyQ4yKteSCjbHYQgdYnPIxec9h15ZLbc1NnWDyW/6Z+UeDkD+ptJooSqqgRtHLj8Be
Leq6XdHWAVikLXhmQeK74rCPA9/uXnvqeaHXuZWZ33pKzOZZVNOCPeAR53HN5lj5lb1K2p7fyflc
Re6loYgeZgEyrPJs/zWpiioFvF9HHcdyzmWNWUhfXBxOvjIhBQ1y4xCaaDCItKuavf/Q/1UNdEiI
Jcywqp70U+BCTpH4Qtq0RM7hE8LN14GTtLMyNm+mCLL3nlDeK98GYYWqFuy4KAX5ptYyeevoGAw1
RAIh3UiIw/8ry+12fAdE1I9vL/J6DL87LdG37ChoDn+8j8ZFEpBIRLEl1LdfH8aQxcW7O9s6FOOr
oGmigROQnAALJhxbB5i6LC/q5S1Y5HDrpkxlXhmCpY0jfbXTznWqDxD94Ndb/JdvuAILZqvO9B3V
fN42wVvUhalBOZ6+oR3M51l+nYTBBwwuLRzwjva2LUXJAhH1qr078DAGLQKStE+hjSu6fT0CZZ9R
F/PKeQXDsuVJTI9fS8yAcvWn8ItvUI6rOhUV5P5z+6k6/mAtGYDMT4N+RIA+00pae5eVlQBItLfQ
SNQSUZXCNkoKXj3Dc/hNIOdve3CbtYc1EsfQArA/Mb/p+5XJj3AgUbeJIW4kR/3FUp+JhTo28742
/cuOLTVHEMrOugMVIidfNV0lhnwmksRod7lwMF5TPu478ObiuvQdwjL+U8G3yFtEi1V4OsolTlsP
41iWHoFAZSmeLCyDi5vCjtIFEra72wAzA7sqJFnS68M9OClZLernKsAwSkTJzw5CCoPrXXA/6u+Y
leBJH99G6JKOlhCnMF1V3fjZvRATY13YLcyFRNsPOUcEPls3eUGGwJQBeoQDr9SdWRqyhFGtCzAU
CJXdVkv4fmI7TR1membpYUXROeRETHnXJyR/PJjL28IcivXNIUbm7r6emM7q0j86RfiZ8Rx5m0FY
W2g8XzpLbDPeFQnAFgAge62GVX6fTsFC0tH9kDAkRF6CDBp7DHEKyD8NgP2ZwLac99lVCJD7lUWe
gO8Zhpt8QiPt7QSvCb3UG2gUu6eAK0eD/kpdv+rgUsK1ZQEmp8T6/pq63/WQ98+BKelvrxy5bgC7
wnIOd43aVeYKYpj7KlyD1Zd+n/Pj2lMwJw4OizOsx2qzCeStrnbwDoxdzoYqaIR9QAWF9CWYBozW
E4yyos3qEvWnREl8sI7njz9+TB0/h8gqh8cax3MYRnoTtECBiMpXnvsT5dszLQYm1YXK7vrC4Dch
3lMSe9P97SWOlGQQR4gYCg/Xuiq9aYapwBvjW/BHn0exGH0RIz3373F9fWsCT8G8ev3KlPR+b/sG
tDEvr35W2WgIKOCJG1sy3LqZ+VuDWQNhVOvJS7n/D5Y8JNMFowWHHK6NQtt2AN29naNVv5v/velS
pujhVSp/v4xJMpmXwExswdK9sbxBu0CU1AAp7RoakEjW+m/fN/oiYXOU8NgNYhpbPkwcVaH8Udoa
ZAZ2Wmcvmb9pyTijjLLJFxjBd1HPDjwsXo0qN4bSaNLA5BCPiicNo8CxAhxhRjBCeTH2W008FLNl
ra8c1Pm7BJi3V7m0ycw45cPu+F3a4DE+IsbLNzqQRZ1a798g8BIqK6PtUxuwrl2EJlGmqcSiENiq
AQ3hQj4sBGszgyG1cN6fgqrJMR2t+qAKDgdhIQCRODVaIQ8LsdTKXGw567N/9CasqDqMrWCAUIhT
mx+r/KuukeJJ2DBi5rCv85VUdZu0ocx6BfkLNqigsQyT9ScExJl7ar1WGnQLxJwcpqhLZe9LIPsG
UP4eXJryXZ6lRtyiQLjfch+dcawTkXKJnSC7DGXTzGLJx9JF+OyNUi166b5Rl0QVvvclUMxurLcp
2j6jXJq57q0iUxDSM+NLlZ6iF9mz7DR9bWHFA0eP8f0KI7Y5S+R44JUJ9uG5eRyV1+lcfujZq5bu
X8DKrrzdGIE2nOaK0+z/uQKrGIhuzIWDSWoHXAbeowhKMlptfY072N6/ze195k2DWUaPlXrum67i
rT/xeEQ+zhT6m78Pj8+ffMN7WGQ6+n9fJB7PpPIyxJPZ+7CxNhYxRTSXHV79SkBujYN72b+riz4b
SLq1rlLbzTKrIK5nOf57q3bLz5Jsh7OxenBDET/rMJ1paYXOzfvgwkNd5woly1KDFt66gR7tR0LX
CDt3reNH2U9TMWRzuxSV6mOjhhKbi/bNEeY4EWakZblOmm8ORLFlBsHls/zgZX0AvEQRRGvQhd0I
9wsMbgu3uMP91fMuJhZ3O8QJwCy0MVZlUg0dCFGbk34eZ8MS4s/++V5y58penYtPDxzSHf/XqUt5
WzEoqsnyvFSVlTsQ3/Jq8hHz0u7EkCuK/bahQ4iY4StvmlI/nKfxImUUkINs5mPZc2jQDFObC1qo
CsftMqfrW8i12gC2c5GVcvO3gyZQtSNDhEHzSgOrTmN5LnNS0EVKowF4uLkd3z+XdBN3FlxlsXsV
acv1Oh4CnrN6Ct5SxJHKyDJtsPtGlS3p9FGB7VhlA1/pejlf+qZRCHcd83CgUFMnz6xHlc9P9RDM
kKatHHxYuY3UCYEIuGKY8R2OA/4l440uiyFJvT9QIsWEYq9y2gEAZ06RS7u6jdNEx+w083SyMYN1
/Dplthcg3rDw0/siXTiQCdyhnOD3fxTQMakTUFWGEABX6LnpYH7lS/eMWVBu0GsbpcV4V1veg/c+
8XMl301OPY9OkMAdeAL6evNd1UBchFj+4uYZkpIaYUX1/ATIu89l46c4hNPF5eWt3s0vfvlCWiTE
pe9urR75WCRHTYs6V4jzy9epHvGpIkVeBIZJRflP1vuAqRDPKXGububIB+Y/uASHjZ6zS0r5CuN5
kBUNV+Udc7VNElApkF1AQQMS54XOVW9qjMZf+ZtWqi5fYscYiOeYoolrdv50/kkucwWff055lNTC
J06QzEI3MVCWi2fCOwm81/TBdgjTNvpT6jKptw7tsrNZKjCFzT+aPjfPAP4107RDkewNkZw1UKA8
3+DVgU2x70lXwCsQ7vVpjDcuoCFtXIy7fqXoP9U0Y73OqHi3hy5fHWm99DjQFUjbldElsSf5RCiP
5CEgi5KB6HjitDoHDprdd36rTaiiil15FXzIcAV0a+VWXiVlcfsl+5/YrIPAPq2IW3H9SxFjFrI9
yLlBqA4q87aAC9hizvuBBACj+jgFW6iLeJ+bc449iRXpRBxkSH6vnu/Smqd5rq7N5DjVVv7/FQM8
8aXKWcSg0BwPzuiwucZ1dSgBJGT8tNtzxDWEFz2JGOuQyiN3U9zgZc/UnqeO1yFHNudW5Xcz/9Al
2dwKvOLTyfRsjeIgTTA3YymeEdSJOy0YtsoIAahezzAXLvZDSECjOFysTXGEcCAnMyNF5lxGxhh9
Y65ZZOThKG/O/KDETnAP5tBst9G2mWB7lPUfLt0cNFtQ0Ym60QeP3D2FeBUyEEHuiEMI5EO+pIZZ
hzN/9xQapvgP+lnYo67Mpx4lik9dbYQpynSg5oGar9VHdDiFksRHk8HtqHXQwzv3uJWcpIpUn/5m
PBjbKMVfWIiJtXrSV1RpE5KQ+yR+R5uwA3dpHFPC7ARUtr+aSnKwW1Jan+E06z8ZspI3yc0Jeqak
f3WQGBk2Q4GlR+QbjX2IM72ZBFhoYi9o/wMdhg0ydrz41Cwb3DIbE27eIIEiDPq3msk8ZV5d7Waf
Jb1Qt5kkVVv/vjybEBZxe6CCCD8Djt7oZuYwZhcLnfnApwuE4bzrSqWkBbXugnFpcNX0hAqIa6xQ
P5+jWuo8fHTwdPnDhbhL/gdsoB5G5lqhaQto9FMYhh9m2plS3So4JDyYgJy1uVXPbzwggWpniAf/
GnFWw/5p0pTj532zG6GK3QDP8kYDDC9J7zZgWdkTgQ86TyaiRkaKetWQkWcunnvqbvwelNC6L4n4
W0pNUyAC7lrrQKVRGphHHKgG1qjyssA2FD8/86rnNoV263ictUbUDIH8Dj5jy9+GptfRPyeNlYuY
6yR5y1MbnznLGJIk0ysNDSzlCp3mBdjecc5JblQaf+OLW0RW2mj0z8d7yqn9nPMEgCanYxJY9W5G
6LSchFVsAQBPNyER61uC+BJvZrBUFyOHXvtbOkgc6tCq0RDKTHMN+ON6f8iIzo7pIY/pXOjN1bLy
MoNp19lTWMOJFAPnMwqjZBNxLGDQh6FyP0qu7zHBzWT4eyyUpo8MTIa+VuO6R9QURDLesrcoam6T
sPXUakViWVupwXs4PKBQpuI9k8TZqDK2KhFQW5NHpbVpPM32GKyUL/Yko4BB3ws/baGCIJmDXUhP
kIw8P9D+RI9ym0A2huDJZdYveMev+r5G5nbExsHCF+bsvkrSnwkuodgSRn+3yFVAIJPYZCuFDGnL
pjxGvEnORGZjltbP+VD+u+VYhj2aQiJx7iM+wnbczHuFSejKv4jNvLBs9ofQsglqOdxBeAvPEw9C
UwlWeEP1RR6QWOaHaUi/s+7NSXDKH6CZTJbLrAHluUxddPlEz7s6I4q9Pc67+ZQkQe0Kx3hTzoDP
qy9x2VxbTF/blvxFGQq9feuUKNkslWB3avd05qqyEPZhCpOihx00O7v5i/9HxwFPmzY9kv/5lxFr
6Gxx3m8K/aK9rJkko8za/vjhATHepGr7TWwclgk+ZGk0etn1jMF+hn0WMaxRI25RQlJOZHN1XMv2
L0nA3Q4SsqkCR2/nOwfn33venZhDdaygHRAH9NFfNhlkaPLTTqywTk+ZltSLewN9HgWJ680xz8PS
t/ynomtrgMp8VYrwiPxOcExrYvUiEp/esDhhlTL0n9VdMXQS8Z6m3fY3unwCkDzF+3TZxc80WX1D
x5G8+SALb+bmJaJt2PmUQAeBTzpQsLwQqj+ws1MoayIZIEu2uQpGS9U9n/RAZZQvry/ORyJShq2w
mPwSxsFxTyJM77hsu6KxFeMN4LB5LDFwbkLow2VJ+ls7usanZcSwW7C7Sg3gaUFbO+4qlybyU/Mp
IAeVfTEbiphLcVwFuY6Oh6CYkDD7GTsmbMSsktkiKisCTC8ncfY/AGhTMK8COqSw1WI1Dr+tVaB5
5GiWLysq94ROXrA+M5I/1Xvu/J+kiTq5TGEMRyRZ+3vgJkPDmx6J4gK0U8pwyB8yjcnDIkPgS6fT
/9CEIwUYmsf5An7cssCoqQriF+ee7r2dnwjUqE+ciN/eSEUmXf3bGLD67cs2dPJUQyufbeCuMa9A
xsGaizglVv0jR0wzCiOjkDXIZjU5FeRerIAVubYw4bRAmINln0qaNBHX/0fTc+ZGNwKujyJruvBY
VyQJZ6dvcCmkxn/cwQf17P3e/Bqh3DNk/0HfjrkjNH3Y3L2I/8jLf5n1Zhap2KmmgxVAdmimTsK5
Ogwga3x7QpsWbaTSXHwJ94yeQD39q/qr9Rf71gIz9r/4Bn/Fz0C7khvuUEXwbzzdlc5xyfbiwars
BolXf8tiv3QLtNI4BNwuvBeKMscMVA5Cml1t7wvJlCWhnNlmJYeSiFXV49RfMtqq2JBBQMv/Hh7G
VIW2QFhl7jg3pqVt4Iz7wfzXG4t8YgzIq/a6jAKqrdbSbL/DzYGFNg/pULQvTj4XPz9h22c0Uttq
rr6Ls7313uSrAF9yEmSGDHTkw5brlieBFgFDSGUmSHWp5KjSexrS8lI9kp6FJJ/TA/KjIAMpkiBa
sR3QANvTtFcIxLppclSClWBRkkZXd6/xHSly5bebwRHSAc3eXOXjYJndCb3yjW75LNWWSF90CPnV
u6oh+JZUKAsOid29AtBraoiguiNw5lCJrp/3/hzkF7sFQRNCW1E2juijIi5EEQ2qHu87WOvBxQAB
5g0dasgrrKSaUpHiGyk343getmMVJDJOkqEQKvqTM9EStzhKqK+mzNHKVnmWNdmiD5WKJMq1EcLq
SFvvHhVS9kDn5VSaSMlzXMUy1AV7gmjmyh/pMMipo0wrHrnt6t89fcnjswM/tKBz1puotcwfh82T
AFc0jue46MVjBCfbgxWCCi9PsR0DQlTN+s1hBoOUrjbxZJKStRZIIIItp5Nf6yAxeqnWg9WrHwZW
bfcXoA0cUYJw3OFykrsvU7j6hx+PbhjUjXvJpJCvIA2ARBrdSri1md3f46bVmfTovUdoiFuW0G3v
nmL4HA/uvZbjBRn6DbwXDf+u1L0npmVQZo2oIdhUdEqLqWCU8vq3nrMDuzCQi60mh0P+aRgiOmEK
EMG6X+x8V/Ti77CxCRCWhJtHxTdoeOZmx8vYdahCQdigpgmidrKxL/0/5XyKI88fNjiL52a+WxOT
CMRkT5Y0I7I0FNIkPMApQBhUTnD3lWfsqw02ot5TqxpIz+LEKAHqkuo9jZCuq1JuwVRidpfqbzLd
Wze+0YCw2tya5KisRHBmhXq0PhfgKtXlkRb4cRgVo0EXiP5AEqR5SI3XNPvBQ6bKeTEEW7ORRvO2
mMrIQo/bxN/emTIj+9CKe9+YI2BuEHrB5Q3nGjhGqMVRjQFmRc1Fi0yHX6EBVUbO/7TFIAv9Vunb
uIdJ3gaJ+0sG1MX2MioL+4sZny4WJSWeHIVRwCSEBN4QhYdGcQancIbv5ffF3ECKMis+NGl6lbpK
F6atu8O9V2NR21vgiv+mA/KAur4P8fFZ6xXCPYFpR0P8gMPevxuryNrMqrMPZ4CSesdJVo0p0HMY
OR/3o4SAp5xSTRmzPjIxTAhvbgbw9fl/L6xrhtD7okB4KB/e20CFptWdM8ulmsyWcgAt/ZoaPjJ9
Q1EaWYWzznEI/ewHnfB1yDfwk74bOxNVyA5kaM88SAob9ZUyUSC369tGhjQ3dGuA0f1WdVAydsx3
zjQAdMXnUjkZ8+zjDxMbDucsKUgYkXCticlotvZ0OwQhLxb7sL4odHXOWp6DkviOH4MZoXaUOJkl
2Y5CswfchzxIRFPSUN0vdnismcBm2o+xSF5pXc1EM4vZlOe86yaT/77C7RcSUdNNe+6+UtpFOv/f
SK6rMRYeCdDUfPAv+g9AfyZ34xi+GIYS8wsBa55zHDUrIntCFPuT49qvwqoJZ6PPg3fS9fi2sNqa
vWoAMtOGIG4RDFWxY4sZozm7DOutrFCdWn70Yn0ElrStHJvOzke5oCm/WmsyUiPSD/AO0dt1W+RJ
VQ4227afSxytosEsVu1INVfD98K9Ib6WOr8ChXGA4NKC7+5o4Olhbl+itfBsRlYVkUURdMlI4TP4
+lBGJqn/nX6J8LX+ZlgJ6Rd7iSieKMF146BOOeFKDdc9NjLdJgIzGQSNob2leaQPP1QLOggolfPw
c3HacBOwbQBTLQhlxe7P46meFSTdUBZAOUXHRUS0H/2MqD6qbfGMsNxuHF5nLJ1tPFWEzcLsQrLC
f5JV58LwrkhbqXzki27LnNvCHlPIepH6+tKqnyh5P+G/tc/GXgObNtjGJ9pA8zlQtWsT/rgphhnS
gwnrfyv9LIx5HWv4CNvu1R9H+yfkWZvPsg9MFIQ73Gc9Gw1gPrD7XeG3QYt6pbCGVuuSoI0elMMg
toRQorT+DEbbpXd7NHxXTGd/EAdhHFELa1Yb2DpFCPSUAseZRolrQk9cPKCfzZu87lvuoYqxnnNG
MhaHd4vJSfEkDmFTz+aGZVjWtI+zEMhpLMrIlI2GiOW1eLFnDjst4RJ2eRRe0vlXwKoiyTSSqLzE
M8OxyYQEvz38zBkarBTOLc2YDL3r2mDdib8k1ZbJO8Ecyj5rsTYnJ1xpZmnXf+kMZ21e8x0DOzKM
EQxVf/CxoMfQS6kdvAmX0maJkk2yE/gwGQoqmJhojMQEacAj3ydmfGs+csBbBmOif2UObz9a1ktk
utTsA8V6mg3ZpUmjo+M0xuJcButpZsGMMNC1mgPxLjUGVQSXcgOKcsxYZkHcvX22AjET3fUxCQlr
KdgZ1eCmnWpry/F2OffqA64Ro4cDn23Hiq8PTDyKHOurZuBG8GflxEr77jvWcEzHaFOVVMLpbpOK
szphJ0/DiR21HGBeXvexU0i/hLUHbMbVsBu8uMHEAhn4NXPdkK6KGPb5KNgPvV2Jg01L+BEsIrxc
ja5GhyAu5IQef86d/kIC42HAJOF+LQ5k4SpanEKEbLg0WlIazhNcgb5XyRhP/G7VvhyI2lmvpBcF
HNqivyQL00MdOCKklK49Lsl6dVIZloNz+jNz0vMRQ87nXVIr5U9RjyoD0XUqTjOpf3RfbxqTuZQD
8Joa2UYv2CgGlgbx/tqvxkTG04nyTD3gjyxfgo+zxQlRwmtpzH8hBY4BOEXMQqikndYEiFRfOiT+
RqOVPeLHWryr3Vu3LBMOZOsvwNca2TOQq9/dUyfrmSLUbcrey/Qnhw6NDhZvhkMlJFOvSeATtej4
+/FwVoV+jpZrGSTuizVv13YvBY0MV2vvUrlVCRJD3b35FSojbTU23lv3MjElOEt1+a24UTWMLGBn
Qd0XwinSJedZw073evPRgd2rWkphIsxaVO7BjGGQ7wjlHOhCc2YpO/vwxWQL/3R5+KGFc/RmPsJU
qRwltSzu5jhe5K6jJyGuqSk749hi7n5eG0Wimcl49dlJwTvzBWBjlHy1py6LdCU8OOHOz1luJAwE
an+usxHtqfhEAHdEm3rlRwiwHc7GazxTEv7kmW38RVMpe09gOYmBqKHZL4aKPTDlKKTDiEDd+c5p
QPc5aBhlWNtGE8YUHssg+qhYgYp5qStQ9/uEdgZMd1ZPeBUKd002qcLfQBHW3WBBjuXSj8qXkCnX
VruqKNDcL1t/V8AY+OD9K1nq5pHrv21JRfzuI5rJhv/tFafpMwVi49VSFqnUfe6OPHAUYw4GFbQe
U5mIjWly2NdpnmpwbDYz9dTfcUAmp2/jkzv9fW62b2d6LlxErh5ghNUFFPuGcYAk6LAPwbL45g3x
VX00/AzlC981Q+BvOzqm4ChIk7lyU2VfHSmYamzMd1eTnqHPkaC6DxdMr9AVt4gAXs9crQF7JTEJ
1T00bTFnx8FUxD1Psuacyfxnym9Gu/oWzZmD6PZdNzOBq1TK4J6cQvNZOXxF8JPrh2lYUlnvgDSr
p6SNwNQFf3Z1s8lCZLr85km67rtZdAQiSuNejCwElcsyAlyoKKcGCQAoN26bCvqmZHZ1wEMoT3Xk
Yg3i3KvPuls9e/6ausg6s2kWwHt828SVY1APscJkSJy3rf80ytEWFBLGHRDhu8U7XSxgfZoyrhLI
7CBYI1YU81/2PsjIklespIUiLZzzmpvJfWfRzhMPNANXeGVB8p3tKvbdVCmesyLuV88ibOYK4lDb
jh1f2UxXrdf01B7Z3DBtm4QQWl+hO6gZnMbT5q8iXKvuURPr1R2HLGe+qoXTY7MO13+GSVuHbm6W
3BATPBlH9A7/j6R26yJwW3VhlfmE6tXnmj/IPNOxrQsQWZMxLSqYHQrdw/X8i4qmcwPurCL/qZrP
Kloe/3XJR3BE4ll46v3MOb4unbs5reIhrwUDLHra+S6bQYKt7FJUoOh0uiABC7t5xR9mTNZAhwZV
r7/1i99Y0kxvjQ2sxtIwlSa/bRLsvjYUROnK+Vs3k4jnUMkM/ZDmfwG9oIjjbxXKMcZzdvKK3+eP
hn1sfo+v/9Misn7gykx1cuosD7Ecg5ZBaD8R2fRwXz5jWG4pG6f8s/hFZ5YkAV1Y0YDBz/klV5U+
TAiGEa1cwaylXjpVMHwXRStga+RWdVS54wF9YUP/2GZXEoGOOhJLIxTFlpi+1H45u7rN6xC6X5Iw
VIKyknU2ZzXAnrPQGqlGe9GuPP+ZoTgbeN0LN1Kf0rOU7Z4c4jtmMSAuJoBK1NNzNmfGa4RAvWKd
bR4q0NmwaWlCLI9RNWuAtAG9dOcP1TZzdGTU3NSGyIn2wCvWIPrdxNQ8YnumT8blzYMMP63W7Psy
dKjxe4M/J7FUOSxAerFuNcYl30IimyCrKxmcRONmKZg7B1Wol50m/Njf5Sw4tHGGZ9FLsYlehtgG
RnoRHqd7AD08UTgql7TfMHgsv367I/H38802mANv+crzBMh84XFGWVM86rT/lxgKUg82dIkkkyjC
L5Nx/xxBeIWUb9GqbWgAP+2Gq0QkUqGvl4CC2tIjfijX//zxBanc3Kj/q/CMPdJxVJetzs5dFNya
eQbNFZsH+Xlc15Wfl3JRZq6t/a9uZRrj+PSARPe9Yh3YQ30ohvPLufgfbKZfLNJOyH/9rt4zyjIA
LkoU2K4dGomK8/lxbeuyTnkmWrvR9M74AENUvh/eDpp2SDbnNZmc5I3zfxof861ttU3WjVwXHySu
nGXdzAKneCVeDmsV0ZZZmdWEGW7xMhxY2mIupgFJ8x61QPIaCrhT9CVv7J+tZr4RwJjeTWxyPjdz
O7i/xcYzUtLX6WCTNL7twQlmr69izALUDGLrpmsGVrl7UoOCJJSsWQUDuGzVP8LaV2ABVk+NWSyw
Vo2Iu3KbiFGAPd2QG9LcSw98IvC4R0i8msNLsa2po2R9Rzs32iO5mOljYkxl2asudIZFIoSeVB/+
K6J4l3z1AvjKvSBZ1P+h4aGI1C952oOOXaR6lAhJy1/9kysd7oUb1rcK5c/PRh8tSpLaLa75/lFm
u70oz1tkDLPfLGxdu9klUCtSt51TIo8FAM3E258hz3nIattqw842KCsuSCAGbA17g+pNasbxNjD6
lszs7pI7ZKJkZOZN6fRdZAgtTJa/+d9m60KtzEtfgS1Gv5THJGcJT6/1iqost6tDPO90TsRlc+vD
rPWgKulyJws2+wBdXeGioQO7GPV3h58NqB4p83xzw0XlpugOYWf7K6h1iX4/hPytA0H+mO1X8dAl
uaeAKe7OejkrgiGQS1E1UGJGpRi0DjN4kMwmeFJH+3AnX5Ttl7HfOhik//1fut3RjQ9yedrg7I26
sADC2Rce2gOXHD07c6bK0AeUMPi/9ZRdW3UvGRM7egytdmuS8+yFVYSEz0el7Y7f2wVXbKuqC3fu
wUImnJkSjmkKWisuOrt70AClRN5eZkjiiGRu6NQXb4+ig5QFN35WiCCdv1wAYtWZw6tymq4h9P7n
mthuQBE8F5aVHJPP4niwr3uuXRlD4QdhmCBJjZxdZxAuDzPNoV1gGv2FXPUuoyc85i31dDVH6ydt
oMNXGWnKEUwGRGOHxJ4GtctkywSqdFsMiFNLVlhyB78UOPz47BnedmlE92pAgEyNaDpd/Bgix41j
NljiuQuQOw+MjY8TfrWv0LXhB5PgdRJruI7stFiaF/6qD8MJXbYAcQ8Ea0Uif8f/SVhJ4LSo7qIJ
YbzE+SF8YBN3V8uvd3Jt0vMoKlkLIUmSH6p7Kkfyy7avqMj2O4uPoj0Ghf5dbgMJpynWdcwA1Cjc
lFBR7t9mewaWGoIfLpan8iFVCO9Y8BBvdVYoBUXbGOY2U2qiqH2ltYV6IhxRVJ5FDBthGeehqrmZ
6RjRAuEuhL2+pji3YjwBQVWnN/Q6wvtIoTfjQ2YXOm+ZMHxURZ1epbJ+LcAPlhrUVZazN1WAbRPw
OWO0RdWT8r92qtZRLq63LcYAz+mwvfFUdP4DKneXa96+zBbJqon/VKzLH5N8IzYOK9YLeVWLLbS1
FgVv3eH1vPEx64MQdQ20M2MgixxhsQZhOOCSznkHDo3g32ogZfMEwejJD6JjbScxTTxVRKUrg15X
aypofCAq6adsGLlw58dUNzZtYLfLyLEz6eTfRR9cuA+mbbLRQXAFCxYy1Jn8D3MkMOcD9r7ZVENu
y0XsKLO1NUQpO8N7YRDKscxTYfVcglvvrqWpmR3FNSheua2CZUZAFeHgaa2+twbLJkopPyLSusYE
EC34qSGPo9jF3OKEYmpuNwZCdgKdH+U1l4HwLHuQsnXyMGkGWTXe+CdwlupuxiOhD6ibNX71eQ65
Jec6nkV3saq/S0NAUn2OzGl8ruQ9SL8WkL1/vjqO4nnpSu53ZXkQczRFP64lzjPa8tGKqGPqVaRb
7/Tc6JjXJ0hHltwPQ634R+yP8Z4o2qBaX5j0fPKUmpWurbavWpL9dut6jFfzdxcfKL0klnTlwAsK
FY6TiaqwHaSEJqbmuZEqLlRZIr8QLvhXvylmkATkGt/CJa8kYmXsRVvpP6m4CvKHJG1ZS6aw/Wyr
Y1ahagMdMdQ+Sc7t5TLrr9sMN3esmRSZ33dXXacDWVOa1Fu1fEH1GnFEYcDQ04Oz0oi766hezwdl
ytQXTB4gHKhWFROlR5Hnv6+oLy5GeZhRAgEIScNJYmyUTpvfAx7DBrBS4F/YZCOVnLaLgIxP9C9K
HCb+NE6RNFdyIGHvTIJW5uh8Ik1EPh1TC5rraqdPMp4J2JzpbBX7woNW3SbRBusn7Td7ByJ0df/H
ffWpJQKQEa4XiYP4kGSnCE6tUpSqWq4CshEdRbLQ59NrdLaFvZxtkLt38Dabn/kWNA5lgea3FpB2
NIE2tf2pXNTLLdDKYKfyVyZ5mZTvVchystPtVmRkk3KtrRGz6OhSOUbOa2rWTN0WxFHAUAcup9bU
rcx8LhRyMRbQpVzXaf/iQkFX7OJAmSW1IJLxpibNbHkMgaWQ4IJMKZGvXAOVG/IDysZzCc3S7bYw
mhEOjp+DZv8YaXXfSyg0XASBW9SxkNLayRQArF7h33A/G7kMzxFeoBXWeST2bKO1SVvgdH/DyMcr
YQxU+L7bAp9KT3dVpszvH8fzdLQPcvT0HNDjAVh+NioJDZ/lEEY7CVquV19FrXGYH6ULg8E2FdAs
a+lX3UhMCNCe1bCo/UlCw0v7DNiMuJmokowMyHexkHUzSkh8gMCkySahVkylztpcDizjyjVKqUmV
WDcP5GRlLqhXVLpugrxRoXQXXbfJiyYRbg/LQsBTbTz2zIrqAtIWqzu/nIW5bYJ4mkv8wI3jflPU
QO3Kxv3AXlVMctfTBXmzOlQOueWvO/x72q7l6qA8tlrg6pv9VMpiOnDo579tUYdkU1JnWGMLYjrS
JOW6NNziY1NDnL9dvQ7H8iys6ivlwYcpB+WBoV8EecbOhodjlXvU9ac8gM9THvBPuCaBjKl2IqyG
zJZl/p2TK2yiLDa17zodUACJoemdL5fFaN0+pNycUP0dwunZLwD48XOIVULDqQI82TXvzgfpsIxh
9ufl2e9bUDYRN/ViKnZch/LlXf/IQ83koQsVPV/L/q01NCeTKF3ptV4oLafSZ2AWwVeCxQxRMtVa
PCWp7Le4p2qIITzcbmUpwihU/8o9GP9cOTU5DxxBrCsGE/K7WgspCWztKTRRInWlntT4iMiSN/ov
lZv2IMhZuUuVMKqB9LaltsKeDFa/vWGpoS/5H7fY4/Z3nEk6sKYc1juEWxfDPig37xVhQhTHI6KG
K9kjeCDCN6JR0hRGOcIrCMemBpuoAKpGpiKuQ52JdFC2DT1U3cG6aH/BMB+CVxQT15e7/0/UpsJI
Mbg+wBE/Fa8SBRj+Uzc0yEaRwFF2s8Uxa4nh4HBZ4e9QuUF7FUsVagLzI5ZlUQnlg+Fpa55RWENN
seIaf4okfR6MvfajGHVPZtWVrn9GiZEL4BOE8UAhkrLvEWVLlOmefJXoKv7KbMygWBRT7sxxlAV3
v2I+g1c/uHBwI5ae/Cq412RoYHbH5/+rnFzKMLZ/sALyLwQIOGdOVQ0AYnat8G/3Hh0zZtPtSmyV
5t/+yyjDtJIMieub3VUvYSr3tBs76IFzhTk73b+MY/zArURYqwcote7Ol7LBLpDu8v3GLFIZ/we+
cFmF6VZ23xYnNBHI2mc6Mq3OGd8xQ9VHvoAvxBBw6aIfWFOKx9NiOsY8dCJLfgSB+YSDH6REUvQV
Va1Hga9D0R3t0roaMikPsgVkCVul0/38F72HwHKzAAJw2Z6YgWlCmga87OCAkcnJMUNrYi8qe60B
wY1flhM5Cfcm4a3DIxf/HWtdavkm6dbyrfc3tmvFVkdcqUJYYDBMCJUfwMKXATXg56tn5AwRPOVl
boydcU/SYJZpPtX6bJPQAonDBo82oGGsO8rK1hOrVyTnZTALnYjH3ywnzj2sXfV9fKFogXsYC3YF
T3kkdPkdtSg9Ld+wEEEwo9iuwseXmXQjXW+2qnCySJsEB9ibEuDk+z/qAn+Ab4rwPzFXIepTAvFj
/q4yWjwhXFFdz+HiqvN32uhPw4NHL927Tcx9wq9bRMgznaZ4RZvNZWvmOTxWY1n8kRM3br33QJYW
Ro/zjhzDczfRRT6GNh0L7q0RLOWf7Q0sG8Mj3C4CVqxPQItIbvIKXZmQ3OxjFbHerlCvAEBf/k2W
oXTcJI19xHONL8mflfaAqxZDyAxQOwoogyJJLcZbhhNXclNn1ZTC4UBmarD1id707oHtobms6MJi
TiV+yIHn8CUx1G4XxUZWZXbzEtDxMapiow39TymObNQxF44wUtBanEhQkFlZ+19Ru6YVIvDbFEDw
CrcqY/+FPYkPTLZPmWJPbzA8143nzLR3HV4ohSxn842T+gFWRgEBaTSjHNm+0UlF+8YFKBj+Hzqj
GtwDRKt5pgRmhBz/jh69pimSB9MDtDUsd9lqB6o5fLUar/33ras85kWav6SACOD3e9Xi+ICluYdx
Fx3iUxd+TM2V7Ku33ls1H2J7v+s9Ja9TLYKt4tla17hge4C74F0d0s9Z6jJ2gSou00P37YUyFUdy
wrM7ARQnyOemQaZuWDT2aNDAxTtSM+gIIV/Qmjdbo83QKB/E5zmrEngP/rCUN6PMLdGMn/8LW9Bf
EMqHJxtCZCDSLSsKFWnsPM6p2GE1UpWlhjEsK77XrORZbJ1mVvg6nuzQVaqYfB2zLbmZG4NhT9oB
oHNVa8i9qsIKcSfU58L7X5VUadDwyxudGi7fi1aInMmHjYizM3xptzHFvKt2M9r0Kdjx8pBUIBYT
rcZ60rh5v/9H1+7tNvvBdjUaKAhJGPeBBOcfHw42JAATXVFSkWhZ1XBh2Lb5c3lzPfgCX6Dz+D3s
yPgkwjJf/Mux4Dx5xzySZKQ3LkG25yKNGZUGiG7wbLoY9dsR03A2Z9B40mMgf+CZyngzD2z/l6Rh
HgZ/jQwyukygte86p+KHTv8kh0bVwSohzWOxpjBfI6+LxMX/fzp42PADRd6jUT+6y7f5kGYIFmDH
HLHwYgMIr2l0lQGJ0lYi5arHlnggg0j2aRdzM0GLlVddMyaFHvGcliT1x/kAjXCekJYDjbZ/XcLK
sNSVTzEzWvdTgTFciWjKhEvKDYfGpkxQan+MSYBwat9hE5Iz7cLEbNMiz6Lc4MkqXCoZ0NRwonos
U4lk2t4gKML/qHzJ0y832ASlLJ7mluBm92wpQ4n65if9v8D25l+ORacaVEnDuJ9jPKVOaBqUcaNy
mOafTRxbNG/BuAE+8Y5RlrIJm8oF2CBFl+fL5ZfqM9J1hTG6gwufV4rer6h0ML3jvIEyvuDMbUtd
ZGuUrtPZL1xj525SSpE8yokqvw/EwYZdQdq50IikW1c5qtGfHq8y5AavTJRL1l1CkizYau3WYBZ8
J+3ofJs9Iy/949WzLYuvU2RnQTbklVxSaZ/4jHxvDmQQciU5YJUTW66rX9zIXSIuGL1W2I8ZghGW
euXZ0ucx4o+VnnS6bZSxkaIGquLRIoV9vAUWEr9uDWIXocCH4Rwdux6SmDd9PaXHZs6F+UGjting
OeZrdvAHhAvbd397OQfl+Yn4xKGmjy4bqaCKpICrE7BQe2cbhFPSBP/E6cvheZA8YLYUHVscgHQ4
Sa3v545fkTWyGsvKUpZ7R+81g7ybC/EyQX38ikvbhStGqSRnAE/ocN/iPgHL41niiDnWQgZwbLId
z41Q2QrnXVv9nGvgR8I6XpkXJxB1pl1wmSdZXz/kpko0TAqW7TP1gUEjBltxE4bGD3hwsMYijgNT
SShfF8UjKS3BZUAeo6E5xo4OvJpTqci268jBBaH6pGGXmX0ciAKhZGRlRrfE5g4xZTgCPiNFFMny
HrWKrfHZmv5sRE9k8+CT+pK5mCkXL+xwfA+mdq/SNYQk8O47hV25r21o75o5U2AiM3YKjkUJ6/5m
hgH+pYRxzKBHd4S/nEon+uGsug7LBSAacoSiWS5GE3LkBC7IbFnyXDy8BfKb1BOjqP8L6EqIzydY
w00ZRE5cNBm9mZb/UX99UfqcoiZBIV2UAX6ozxQJrLuGH88IYbFBP6eLN9Bn9ji3VQ9yNCprI1SS
aWNgM/jGy2JX+lGBRRU9SQi0iSy8d1ec902rZjwrzdvg6DtW1e6Ma3RUwn6gM6A8pLWInNklzyaW
qrKVZIHEg0lVnxVaQR1AAt6ndGmooHOEobYr17HcCZarWOM4X/4uNM+sO9nOWg11NdgZrj45N6lp
TWPAWIMJbNWkd1hL6PdfROarS4tGSAu9EhT8QOAuoa798wGrGo6DxdAFjweXMw19NTuQYfoiVsvA
im+gU06TIEEinJgYvLCHeStX1XoR8WyEKIPrcmKfhCRDqbXVj6uVBcdW+4DksbCY/ZLT5XeXMI4R
nPR6g8RtbePor9hZKzjmuiKvxjrNoGRmvzibNwoc70YTUTVwRuuClbtX/ZLhXwSOYTKNc4AmmOTj
cIbBHmJmxTWJ0ygZGd5Cx2lGoN7nJh4RVhD1UDCuDAWM3BJLY2PeRMIuYkcnGB0tTMSvUY4ZcWph
OSxPhnxXL95qi/eUnQYaaYnm4F0fNdHwfP3zVQ3LDMx4Xu7yzCPzE0uXLN06yyD76L71UF5NclBa
+Xwk2sPcmMXflEuKLYR31xU9MfsPuYVTEJNdB3ivWFNqwRYrJrGQvn3oF3kvYJjO1KBbRyYDf/kh
FQpBeSD3GXWAvQ7hQUORf/DwppyF/5G4GV/bq1xrHsyJPRq79Pe8AQ8Td6LwIVdNGvr+ncZEUuqo
G66kqbbeUDHfGWJgtDi/A452MTzlVpJOxugCo9XONOq5eAq/vVCJdR6If9f7lq6xD9CXzFfLdH02
F2ARMhQ0wBxsQxV4jifoPqvRLb2Q0AGV0tSTteVFlVRSUKdYFXqRUIg7MjpQiEA43Sj44SRfsZV0
qrC/rCE02lYYtjjWOlWzqYARreFMR2KvudwP3vQMdHDY/JgY64H0Q4OgFinZoakMhvfGnOBB3sab
fu8BuMKUTl+o+wCXdT0giAHOpDRtsdE5JqfZflMwEZwPz1+aCCY4GQzkW8+iJwIpgjatuQvNMMqs
Nk8PxPlsms+RowYrdUys6pmXScSMJlERM30ggrP1z7ucU6Bgf8bYfcB8On+N5Gii4BA9u+bpOzEp
aaM7OzEn47afqLH924IglKI78tqj0MZ0hwqXHjkhU094k7RYZkzA/qaS5EbyGp4tR1kMDhRQ1xPk
qABVd31ySN9YjMFP/YY7PpRVW+mPoRl0Q4psUP91zWaTkq5Zsq07ZH7IVW62dYevIel+MDb2gABv
f8iLSX2xkZrl2lvK0ZxAS3OLFoBr3manZqiXXgmT5TPF55M3vfRx5x0qGMEB8gzc84R+LhvgKLUi
raJHmw/L6M+UWrRw1WK/bHe0yz3IAfVqsqQJpyydHPtgFHZZKoHIQSq+h4BLviIg0uEcX1RhqA0K
C1d38iCH5OoJyz49sqAj1jh3Qyhodge7zj7FMNKQ76RXI0fvpYUmBWnjD5vZ4O8H9vsC7k2brirS
V0E/NPaRnAPtMKriLumMDrLjMfp1eO74xryTI73dctoa7MgW9/cf+EcrzwfTMSU2GrufJngl4SGg
gWH91VFAQMwhMXUugc5LUMRqzZ+YseEy2ZEzhl8vIM55CiOq1d+mF2YLcXKvsSVu4zywGCvMuMP8
FeL/SiLm89vXvD4D37lXvo5bl1DZZWDT5z9/vDZLGULpN1LvLDgJ+RTPLm3hyIWCXW52jsX7NLQA
R8nWC6Z/hfViT425Le8ttR74CR0zNFMLSbqMQCoSTdX0R1wl91SWiqDPpmbhvdgM+/AONlpYj4Yf
D29S3v4CRTw/3/RBZK9V4dUEolPz/10GOAuf54sIZGYtmZpzRLIpUYjznNJhneeYgumNW0nLpOQ6
yIg3e4iKTkaoyJAAP4i5PKx5E3gTVqUjGXaT+spLmsLD827LGHFxNmhFUEjLJokJCbrX1Zg/o+lH
eK5HmGvwXcrVY0KpoVh2O/IovFQmWVZjYGEaYCTZGdPfXGoDQViLIia31f3tHq8aWfCLGLgdaBv6
cWVKrFSJ24yMWncYe3oU/R6Psf/d/NMbx70Cna0nnImuGhnXSaeYD/YetjiN9Igjp+/yOH8Jnf0u
LPAoI2zScrHf3QPCPVcCpEZ+tnBpa9zIqmYsg68/KNOTVUtDSSsqeHN3w4AvfqxzGEkTpJ2AVXbk
5scPTnsHmd23Biv5fSpwm4q4so4/JamPWMwzaLxUhihamAgI8oO2J38NtrHnbmZUazncpWv0FZgm
vPsCB8Mb2QELjHodc7bmRVHv6pMpyMTduV+8QX7x1vNH+9l9HgZDaYBu5skN8SD+txp8YWp+QUUX
wTREgwCoAgnAeRPLmLbKU3YTtA55aCaIe5D/pcUQGETqPKbiWfdSL8074OV/6WuUeBOYsbBuBMdM
IzJjy2oFfQd1IkeWT8rHW4zz0XfDu7bDbrZj51ByWKOiB+09izZJL7Zi4l6/788hK5YqoMN11oNf
6blZbW6eRi00wWLgQeznZYrx2L8XvJwYWeiXs/3GuSBZ7hl9HTX+UESkYn71tY5piV8+T6SaJWr6
8r3shgUDp3NZ2vv/liNWyLyN1MBNjyqIC58dEPwtXuAolbwfNU+B0s4BpzQhrtYa4AMCaZPF/3mV
37xeHPUG4y7WnhIPo6mCN+i6B99KYtNCKB4yAShp4TQwYU01erUI2g2tEv5Jd10jNhyu/jESxYW8
6GH7pr7ddCdT690R0t+gZnxjGx+TAGPQmfhaaE47ArXZ0jEMyYUSLbiZ/5GZsmrBBkSVBECxqZXE
EwZUEB3dYrJ/EKzQMF2C/txYofN2zfopiNp/I9WroXdsnKenADG2L0XCa+KKdgsl73pA6+UhkYkT
kbkqHDzDRtSdgE5lX6iXw3iJwkx84Gbw3ck4LNt68cd4mcBKBRqTQ/E5zCZCaRSzqcmO7vkjunSA
VjkcehfZ6m7f4mIgk1XwHmzKLoEZxMYd78d6CJEBDIJFTHY/QP3XzDWJrukd/aljIlpZJkBSqceW
/xO/45CwoG0+kmjLdy/MWI5mocDd0335TXaFEG5g9Oe0KjRUGOmuaNcmvXcr/IV1rq0OLipXxM71
N6SYiWYBaAu1j0Z8ldBYQjxlauJPkWfeUtFyjrdA6UYJ3Yf8ibPR7SGvA5iVru4/5i+LtTmqhSV1
zRk0aZ3BzwQ0FtOJSvmkhz4gGuZDDEX7IL2Aznt24oCLe6cUvbhg+7ItTvaaeM7bGVzPIHUWJhlG
iZFMwE9SPPV7iAFBFZBhQDqMDcX/+1qgzjU3ZRodDBpsJxrJqSA3aiFifAnPY/RY1vPyIruzpRu9
EgPyj6t9+jYA2Fb1Dzt69x9tZYyUVnru2qPn378Yt2rZ7kRYsi5gn0efuL4nDURam+/iTYhggMkN
yfCPAgCq5sa45vJmOVnMgDLrX1V2bBPmb1d/PcL7H2oOpKZ04V41GbVjw+TeBBfvwVJ1TanvKED8
mXDjkDu095TaOtqpIhhMQncSgnymyE4K8hl92I3BLse0VBF+UsZGq6DX3jAQV0QN9r7H+HyfEIrE
gbUp8MDwFOTT1AuYUH2lwb22zCLq5AQoWxehyrw4n7695UWJzWemazXcVuxLGXimsxhhi5U6sQQV
l3A4lUMMUqcuDjYsgxPgueCzRQ55IP8xQisbJiRXsXWkKUK/4qgqqSGq45Nu0voXjgzpbVhHb+gw
yIhVC1mK8c5ORjINlmpfF0diiJnMbQNxuZYamui1iYAHm8sVv/Z71IvnDrbOjrB1kCTTLHOxlEo5
T+qm0qBT301TWL9KndU3ovtIqekgjYndiFjm5wIB/ajXAwNEe5KB2UIbHpdc2Tg5JV0EpcHZSLYT
TiyY/QmWjcNi+5e+GwWZZNRv8WiB4poxnlqWCkyVx/9R/+HqEw4QpwWrtFyFNrEoTWkUcDN3V60c
8YK+Egdrt9Yh83+hWN2B+E5Tyn9YNA5Q00nAh8YtroEJZFk6aVVpxK5YLhkj3RhMxLzNL/2YMlE6
cHaDzLgXnOn8MHyPjXwpC+8W9qPQYor4AlIyam7+CfkCUPGTnYni1yY3cOxMKoEHyUG4Ap/B1JQn
D/+ebVJol48SZb4fgVAfGHBONoSW9mKZJFVTORu9ZsPYsKgKOUA8VwLsUdIExAtcjUiMnD85re7u
WF27xBVx6tb/7nYy7z5EMs8CriYnF/Oml1wbsfvniJWN4PW8GDGpM82Fe8zmX0ocS7jt/9yTsZvM
wZaH7/+By2U3vcQQK9Q0zxR9NMkrb6WPiCq02Pn1tBON0NdJ0ASwr9DTSEr77RtG4N2sKnqBCqnw
mkR+EwMmPtc0PgMvV/pirSesLBOYR5oDHE2gyAEXZRdnzPENaFSUOWSQQrGT/h5yDWg054Od81yd
Qi5aR03b7zQ+0Qau4VJuulpbmT8LkaGMOs692cKnmbP/LKFkrIPEADBkxXpGCj23DjNzr6fHn/Fc
mytHq94obJIPuP7yYqaImPB7tNDthtrawvEIxUW99T81Cl+c/38Rble8hQY9w6z/1ZbBY8dlUf3q
3IwCilIDHryzwJYZYax4nImHyYj2j1Td8JG0RiEgb8y/meKpFrqnCK60WHWD2+qTTVsTtc33St6V
FVZAiRctcdC1q4WBvGa6Ey08JwGD8jlw6uTACsXOKrctnS5F3KgipHNQh7eD1bZU6ySewTfNfKdx
HnDzszgRFnEagXafLlrfyfImIM7Pao9hl2b0zJ5sp110wekD+r6UKtaw5DukXx5QWXGeSFnptN4O
DGafMeu0NKVqAfeUu1gclbOQT/oc10HJok++8rUvT4Uy6sHLbQlSgW97uFp6sKMFXLCe8f+/HbcA
Wys7/EDVGjMYsjQJ6xqLEjtqmfTv1dUzja2L1sMPt4l+KbMVyPIqFRqacLB3mHXtP4SWzJjaKbhv
cf8MZ2GN8l3CXOEj9nto5S77MzXF2UE4Pqo8Y8XTuVX6kgz8N19nqWMrQuGKqnWTkPawd7Ta1cAw
wky4Moqvo0G3u8WtSsgmpLRbzCo0dFcMiyHyHt0VsDzCwfYJkQiXpgTaYXgB5hg85ji1mr7kXkEP
Xx7oCpigtgMX1jShgo4SupEdVEAIhaYeKVSKH87+iFQvs6Q+qrLRX7EqhExPgrslnUdKXcGX8iS5
Ax/yMu5WJ1rSEhMNBL+Fh+wSWQeFdasyZc0wDbCYNgcRDSavWWRM3T1o3FMiunaM89e7OSeAjc28
sg/Dnq5ZTUe9r0q05GZNIlxXVPdpkOhWJ7u8rLF9SHNx+6cgFoR+hq+8LtaVL4GJpMbSCPNEKESo
BtpXJqFvqO+z51WbdqgQDlfIa5XiqCH8rTjahbGKwwmhBc1OYEnDnddqFQBuPHOYnLJ364qWqICm
LFa1izscY31RqS89IJjd/IjWHBRwRVeafgno1itLFaSxLk2k2ILIMNAz/Gb1iEj6Oeoh/B3HOEwH
h6Yl+ISic/PdtF9t7Z9BmZ8l4IKt9Eh46bovlLTUhU5NNxnT1wuSKpLGQQd+cdewCSM65uFsMHj3
69EVIhZ6/0f4jbD1LYJCZmWdd3V4GXe6jseGqOTY05Ajd7XJwC16hWi1BXlQ3jWuIlqzcFS5xdA+
PIuA6rTUCH3B3vPMrqgkCE7zEA8i/DNOQwpxcCFksrD9ujSuhbVvemGHHAIv2Hsxqc1xAAjrpH4Q
1h10sW7vtJsVkkNpEiwJ8ljFyOBboYbg0f2Ug+hXyvoSqwu1WcsfJ3O0nBKRzmTnWCqalJB/+7Yp
Ze4zsyULuw9eWNyqzYub8hngRdkplDMRWiOEKXf9x+Xd8McIBB9NdmuN1YiZtPR9l7ZamZrq7pD5
t5dD/Gs/R0OZ76B8JB/yzEecU3OLPSEHg22KlKYQVTvazBjqKLZnr/J/12Q4bcLXVyDFiJvABGfS
2qX2wbwTJi/yuy6NeRm5sex0F0SvZSQIiiJqeE+drNM920r6YTZVvdkTwl+xNVUTLJ+SfByIe0OC
ECsKl3RgunW328tGfyeTxfMEv5BXow9BudTVSvFggm4vs6xtAKjcDodVtegUI3BoPwyzbrDG3yDg
v8tKwLVA2aVzD3c+HVlvu0bxXbprIKJ/2vbU+I55fzG06m9Laqch188cwtZavUGe9jjmVrn/JguH
jftIlR8vsLMZjZ6w/04GiUAh67nQw+XgVrUHDGQDyXekH1p6eL6qLWpJppsfCS+Zeoz9/KiPMANj
5tKNbyPoWuviYr+FyA8+K52INcvcK4l2FN/HCXQvJ0nXirqDaffcUavvLKJu9jZ1T/R6XfqcSURw
OZ8lBhMoei3l7Yjm1L/2zQR+X/KAnC8aEUwzz9pooWxRyE7vnbQOmTazxnhqm28+QsWcUrPlNxUE
mEPBsaGfo8biAxjf1LQkwQJcv7uRFUd5qzu+iKx9QTgto1tKrd7Orv2l4qNdnX40pyBlbaVOnnK+
BH2KmoHC7shTkBPYBbztdqeRdsfxETF5GL2p0hXxBM846CE3ibIGbS845hEiscQE4AA3j88drO72
AZVUwfButnyoOd4J4UL5g2oOT45LQHosBDkpkKoEFm0XrCKxXCXmf3z8xJYVdLEhhkwo11Z/qwuT
6+x3afWqF/gm8SR7Y3nTf+KZ3nB55RGpGnneC9539kwOunVQu5YWvJN1kTE7zRWIAdwCWYl2JYCq
YvP/wEebyMA6vCK1igcrf9e/GxaQNob/ZVsR0d20juMsxDBGRHxDMKVcHla6WeBQY1FSHdr+kYQa
6jDyp+SPeDw/4tfwOtYfZ8ZBMkgcKTENF4+EQ6XTuZB6WJRCIrfJ+hdudIju+iqzwO0hM0NJ/q2O
e3TmnT/tZfkx0x4X30X+7MmOHZoBM5UhtBW65WX6YxLBHXpGFP5ZP/IpMpGZNT4Yb8wjTKv+AVGX
1qp6CU23NKfvJ1wBf2ifMG5Q35PwUHzOMZoI9oWaK9sQvveX+RJhMrN98imhjYPcFziZRUJ/gJa7
pNzxxfAQg+zEQARN4W3UI8OxUpqBbnlxxvBrg0pUx7ildX7XCQH8yBw8tgi6PaBq0RNtWlqz4ebT
RIWkvhIkfM18jPbKKNFBo9HOpG08JroUfdCBjrBcIze4aYPvxksmoKaS6XbuhXyf4JQqE0FHgUB6
TgZ37XHF6TTLQUhzvq7JVu8T89DU+fEadLotXxsC8WRAohsCDyPEN8TpaNRQJGUx1VYgmsuBPpnR
wDSd9HyhP2tPQous89xR95boIx2nqujv5zHlpGTIDnmWRH/724YWpgKQnWNsDxogUvl7sPcDWZz1
9YLQsJ3Ar4TScaE2GBJakccOr2jYKe8fJMpJSU8VNBViVE/ta0KqVD0sa8EW6rMJbXb3LweB+trq
MbFaYXpOMy8jd92PSvT7vwDEmS/qAZAJf1VW6zRAW35HX3xM9BPsx1/XtRgjOGpULL+DlBMM1rCw
tiVRwo92i7ar5Pxaf395c8Ra5BE5pnBkS45IpdUikFlYpXoNpViCq4OWK+bff8Fi66qmDllegXq4
+UiM+kAyccwFbCWMqIrmm4GwC1/qPB4bT0IRzYJx1ynrPzweDPFydIP2bW29Wy+7fOfPqGQw38EX
k9vZV3KtnmuliWW5yDoVWu9AYETI3+/4AUsthBw3Mnzc3NfPTCsvcScuc52qtxSz0H7raNCPSrue
oCo/gHqbTeFLoqaW2poF6DE9Pstr2AtRpiJq7CZc69kjK/Js9IOGaVx5capdm6A28AMJKyshu91k
qvBEoExLEvnUgLnsllUewxJoHj9KfRqnPGDSJ+ZaGUeTdCtdiPW+NCrcVp3W4kvcdAOypYyZQYxw
FAzClEwrm5Qukp9dH3+IDVcEHFgmm0Ms+YKFfQA4rVj5/UisYT3QtAeE790CCFVuLbXQ96UhkI4W
o3Q1+WlGQLWOhH+0zdEQymTHB7k0ffDL0jTjKTuVH4bwvEjZytzFKI2iHfA+mqul0r0wmLlhiAop
2OYqPLTxFa/8FlI5bweI5kou4XXcX6gHmsQ/lsn3BBrSTQ/15TiYHKj/PZNgfDkHtMbzgTFfgBd0
RZTuuvodTY2LyN/gPjzjoCWJyyd1Jta7FfBkruvkwEbQG8ktJaoVllhiaAb0XAaT5b+DXntVyz7u
cn/SppgPIvTPpHvNZubixpsySUB9lOLC8bEao55dkemlANH4Zh90zp9PvIRr4jX/8PnJo7+uAB5b
wsxCm/BtNfG8JBMMRkyoawph2oNroQxaSCSdwL6A6lxDwBN73+OJuRYbivZOKp30Q5mmqhYpCEQK
zb5Z0C9HEkjNv60mJPNa4cxC+iRNb0ZFWksb7A4jTx+w9OzSyyGawYTaEy0UzFBD7qMG3H4CjSx6
4J8DuDFcKH3CNdCT8W3kGQfphOr/oHXDyMk+cMCgeOGVYktx2Ckj3wfmGZonjMSNc2DI0MBNNMZu
SHuy0WPRe16/O0/THLAjTWxblhIxvtwDecidDZ6JK6HMia7NY6AjO+8bltBmN0+2RlkufVknAjYX
cm7BQg02RHlsqo8FjyNdtz7k+YM2WNO6HtTlQWsVF7JwdUWK2a2181A2NYmRmWeBOnHnAhheTK0B
0Xq7gfQiPmw/oIVqTlJBrOGhHRccB3W2qWPnlOzM5c4TApiLKolv7kmR1EF9b8pGSwk+o/p8ebCo
C0CVs21+08htcYyTOsYKHB0zM6nYODtmRQ1WsKpoXtxK5vOPFMsQjO0LJgcC+Z3z/XN5dovD8rPy
buOCzpGd7ih0pna0XCHIxamDv7BDUX3o33fnkksjxDh2ZZ4k3Bws/AYFB5yv9lH8OOoR2MLz+Fe8
ls+zciAbz28xXg9oMbnScb1GJEhrFmIfR5Byvc2wsOqVeORI75ABSygLR3kGGA1as8lLt77A/tjD
1ddUG8Fewje1Ytnv9r5udTmtSXyPlPsBza0InO/E7p0YH/11my/10pGTQ2oyXAqUFRauNIslKklA
QfWJLMqKMe0NdV5T0wcmamgpGixMQVqqDP22Pz4CmIvvlaTiAUUIGYICN6NKV/wYGixQdqVJpsqP
Kda2dRt4QftDzI17Q5FS9temEQHgxdNeH1E8s5Q4WXUANnjXzcb2Wqkgh4KSODwIS+8ZYBE0l6TV
3jiewg1gswdHTC7azf597zR5TQFS4MbJmI16y2ZZyKLyVLMXlRwgnxSOzTGNZ8yYDu8W92PEa90C
IDMFJIsMaKfFxZiCg0VjgDJmo+86pWaFFHppuPx892hop+GnAPWVpqajKPiuJc6LYNN/bmexizin
ePNKcA2PgrP4a/kVuM1XGA73cmrBhvcyRcMImvQlAaSjC56DvesEE7pMra/ewTISJ/fY4t3gVHAW
To2u6nRDts3KLLi6Tcj1T01+spFonpqny8a56Z7sTwiYEFFQBxJUmoU1ZWAeCjUrODv+1MwMolGZ
3L3T/Y7yYTqyO4hg2Q1ELVUPZlmBTUPiZWlh9o/B15QL69nbDKAYDhA1e32AfxT+R8A9pyBnC2g3
RmIjxP3H+Eqy0gzqLM9fRb+DtQx1Me3XuuC6/ra78aPOJHYUbmLcfoCggnSiAiNRb2mmp4iwNsR2
Wt7zPC+6KEfSa85dgxrNJ9D07UYLcdWt8XyCKHjZN6rm1Z+Yr5g6OEEUnS9foTo1zYykkMWdKfdh
D+4sVOZoBXOrm1PDmle80IBQHM9fvl06eCsWJV8PunXGLihDHAf77iXJQ9KupYC6gTGqoPjU9H9e
6AODBjOxWtRcu17EBlHwXCWTZqgNYNPQu1nnyBPxdZycVBce9ZPlFXYyaBsq9xjULoeJ1Y4QvXzJ
9c27K+7ypTm6i27491Vh+tUzAwbYoNcsQy8i8+lqhC7NfSKxEippO6DkBALfD3LI3+SCWoqyCjXK
B/LnA1+Jx9kuzPAMISfKbfJlWFWXmBKW7ZIMgw2gAM7bOJsQ5qEYAsA09j/HU+0RIHtmToHccOki
p2ltMji+Ge3N8JA/OiGoeHiI1hUKnO3dLff1IhDP24k2iuSHXPqYm0ORWHSw0rY4ZvRpzcQJHA62
rEBDJdlF5wzidA6mg58RDjXlAQNODajwY1UqVcKKBqLCsmvytesaH7UEgrO7kIRaaanrsqlJWvNE
tm4R8RE3eO80QS9aDLrmAgs3p8g3R6na1eCBPhzRxZsGi0/g/zXuaFxo48AiTlUS1j4r5g+yiRqW
ejoW7tKfNzOPbdHMxdyxD38hOU7wf5vkayYIN62GVQpQotS7KrJWMwE5Ol0URpAuq1KgpI0Ib3PX
5D1I/43MBhkO+XGZrFUHCxo5HnruBBwPLKzXdOcpo+DiOD8B6WxAFlj1LjdJ9mAMlgQQZybzTQef
HFR0q7PH7NA4sIbCfA3osDkR8SL3DeYoSpf2ih5TM6TazFaMwd1oIC2pI/nZc/LQRZjVseWyTAdt
Wi3o5/rw+LmbVxF2qR7djaElCAS4NydVQ4Vs390yqpFWnQjK54EJmaTEVfJ6jN64xrnJbjB1EgIw
p2gLH4MsU5iAR2ASwxACXM8FgWrxobJHMHZ8Pb7P/Ed7wZI8FG4zqWfn1x6mxkRYh+rZMFcPnK9u
RSa7QFNw+6oZqNKCtdYzxCWYk+sk38nRM3Cic+tLc4/zhd602ni/CuT+FE771e6fmGaN39MZFSsg
VOVS9/P+MOyyyjTql6Sv5AK++/k7Fnv6DbrZyVec7NtTZU54LbXcthpN9J2FqKP1Z5Q5LVTKlRCd
g7QRjJ7RdY+Kn5lYmD6iNVilS8VOBrS1d6zDwWXMAV+bhWQie00JubYWzqRn2nQfQuvMEMQhk/rr
L90MMpwgtrHufzYRmlVKrBYtv9FIIVNz/mbSvwjfL5UDyvGErT/8Q1LBD5Ro6VVNGJasxfSLWfPn
bJaxkAr5ZWsskFqtnG61L0pEVewH8Yfxb1ALpq4eW0qKNy1HtiF55cwf9WlKjeviJ08fNtex+4ii
+0AqqIC7WDwH7N1TM3aKnNkHj1eNQgdcFNrAMOlAorefAJoUTBKQDGMZ5NZLnLwa2U1p3Z/dX/on
k58wQSnpADrcXhPx/OiZNDPs9UAaeJyKmXB7RHCrKOs9l59KqifADPGgK+9ZMtwvMxdRfviONG/Y
xJLHGJx8mj8tkunNBly2KGodTEYTmEtxcswQqW6O2ueqFFJQXpoa0PjYKI/YE+ZSbUeAS3n1JEaJ
mlh/yBt2nPWiAIeepeKMs7ec4Ggm9c2wUCdPgZ6jznCrbgaUkBMgh4w8prbcDXmbeX+rUQ+Z2eZ8
Zz7cf9SfwjZ5ZYg1T6J9s9GuTsCDZhQpsyW1UQipic5ok5VZG8TuIUvyP/VnIlpFr0xQe7paK0Jf
VulymiXXpml6e0BJLJQOw5dklXz53SJ7wJp68iPJXBR09JZDFrus2QQCkEZgfEOh5l8Nzce+33Wi
RWCDiwAFfkB/ts6P6X+ReNhxSfaf2zh3ifNTNo8iAGjFByOz8tL2khecLhPnhVhxXnd/B/ESrv7q
LuZnaanLzCc+5CHewAEMCcqQSlvDU6lgJipn63hF62Q8s8Z79R4ibnOLJMynnKGeMbwRheLgQN1y
+4YRqitWaJZteNCXsTffSi92XOhcuQpaQ5NHa+jcNSxgXVhkLPSNM3DAQrVIDIZ7PMcdAMZCcJdQ
950Pu8eT45V4lGfg1dm4rjYJ3DbDO6SLOBXKApai/ykZS4NjF4UoPTzHETK72swMj49sW2WDwOEj
kXqWKPDxOH5onG5GFL+izt04+h6QEBEi2QO10Aikc7PRuNoxUfjp9luNlRbloQ5Pm65TU/QXGTr2
pgjh6spDx/7TmjiJRwsM2OfNPe9iXtAIWnmob3UewsWp+T1SvVrEXCBrl8NLFpGAE45HiDiSZOYQ
aC3xCKxxyLLkEhweP7iQVnFqBi7LGB2/+QKOPqPumjJ/4V+9MEbl3iqtZxva1Lw+TkkaJRVCM3b4
hx6lorXQ+MQnM8+5v/RrgUNwZ2TvVxxXsiAdAtHMrivGpp5fyO9g+63oUy9kJq0wl53jgx+v47Uu
Fe+VTVj/EQGW4nqgjRtgkU/tcpZljA1RcWnNAT9qfF4mwvJwYrIpfh5CdupBVU86ws8AMHWbZd9+
H7PGXbWyyxPD+r0xBY2FXI4ywwroFEzOz/XLtb5nOSBZWXphDmtU6GcvjJMvMimjuCYjGk1lI0HX
vkDDSwss69He3q0NSCH75zZuOnWlBZ+HsmwqbPfvOBGJhgGWpUf5nVYnB5pO81Zy4DH8L6E+1n64
qLX8UOzxU9hbWwGxXuLRi/zK+Av6GU3Spy+0eurf+Uzj2E4+k4In4xD6Pnn2jtdlE0yHWGW719pE
0CWcNMxHq8VZ80Dku6+ZRmEZxjSyoLjLWaIK+6rxkqi9LDDN61W38yUfJJwjcQppK3ADDo6azoo9
IrDkuBUXCfyg/lk/9hrb7wGExvQiMFk+nqGoCBk7hGB8LpvGyktlfxQ+r0HeDQSlLLtPje/1Irf7
8ncucP1TLZivMxWU/tpA0LBD2Aq5DlMyy5IRFp95Jdt/KgEkAYBWaaLmKmlMNv5mxmtki7oXKF3Y
+9sOJIkuH5VaN9LNGsHKxf2Y14gJrFEMyYa47zXvQkjcFC11coc7+trLDiBVS78kVK2UAdfFrb+f
lapG2iRp/BahvnCEMTHZB0Os+hyjYStZJdf5dP3OMlhVf/hRA96l1yqMCUumMMtXvHUXHAMDNd6E
E/g3S1a56xegcTSw8RDERU29bl7CpjDNMHyUI8HZ97DzmCPw2PUU3C6NEALoRJnzt+CHOIjMr+bx
zF6b+8sFIqrCDk1GTVE0x6BQYTcILKs+PENj3tbS9gnM2KI6oBbOjsTWVwqgpT5lMCMClfzNcWQl
F2MndBX8bjEEL8Ux3qRESrl0CO/i1HxTllIjFTWIqC8DcqekeFWCGrVOuwqDueVBVyRFBLRL/LQm
jFdrgKES5mhVeyOkFeTvUOSddulJ29NREZvfZTgsrJ2U8E5Aewdwtt7SpEB3NSwYYOP8UjES3kXe
L7M5eKP4ZhjxWrooEOwG8tk5J6ANeclPBOA4CkfdrA5Np2dqhNWJ1s7ShCbZ2UB1Os8Otj27gbt3
TMf6JuI3UXNzhKfb86e1HtztrWmG9gXuIDoEi88/V+JudDwjAI0ycZgnwNv89xxFdsDUqt211rTz
kZvXKQvsxSHvAgCK0VjsI52pBOOPh5wnrSsff+h+EQ9uFpr7Y2vwv32+VGg9noB8JpGzNJQ7bRl5
1le2MnBx3qVK12k6ODnsYX6XCEGmgedA2yjvvkhQ7g68bQJhfYc5HQRW4L7OTIariQKNaTroLIvv
HGucT3VwqeTPfRMhfLeJuDwqqDIFdkCLgv7LpUURz724JbtG2mVhUYVkOaWAsyvUMAcl0FTLhWDO
SbW/FWB/GN5QR8c4YobkTGahvvE88l5G97wzGBCOps7jiwObWEvk5Zkyoj/3Zw+qhnO1QmZO5Hy1
zHZKzlvtinCj2a3TXLfmeXW1v2CBy2AebMw0H/x+h1Yf/dinOCKby5ZbTy51v3vdnS7ZTCN/c7TH
j0ec+CHQW4a39DI8Q/LGBAr7K6d7r7Sk4fzyZRWYkkTHDHRlkzU0+JIdm5ygzoOKTC7EmtZK7Wgk
imzdQGXxoO//KQxezyPRHx0QRB38TTGnpgyV+w8lIxq9C5a1EaD+n2rZF+2MgZURSbhHKTwlV5GM
uMuc2kT9RfxJIVCP41SGdRutd00QSk6PPs6hc4pFvBPJcuB2jG7gG4i9XEXSgy1ku56D21bgzMXb
iNflkgwHnMGzGflu4WC5wNi8LhNnpDEZgSE8TuUi95wlQ39/oZo24deYHfTdQrmxbBTfnw3XxZq4
NtFSTgoqnzjVLWGyo+nQj8lj/hxF0adHmC3RiKjI+hEfkquGMb9tPWIBD46wOPADkVYLEf6xSqOn
Adca3izMtUPu2gOgCvf1eYGYgaEPyV709+nxeoaQeQ4+Biagkn9U7KfjohHKMlhmUR3x+3yb2/He
+924CETFQKz5f/pVNNymSjT5912kg/c1wo6iZuXFQVlWXqy/Lv+x9fa/19xF2BD3GaEWNyQ3KRXu
Vt07PGrWhFgfmTBvDrHEoQuovbE0vIQitjZKT1HYDASrolYvPEm7YTKpQ8IbB5Ro/lBH1h2weCpf
5T+bQ2EXTbTiCwOH7hXMEyOv68scqoPfE4sLS2Dl/luALdFY8AeVk4kOJO5Bi939JotXc2xXq2T7
9KZ7b7vVb8linvivG2RhMlnih8y7hJbNOG5dsCNuZCXS9E3zEVXna4vrZkXL/ldoq4Tk2lm6DCjf
dxXnqCiMUAEGhh5mAbbFMlFerq1jj09aC9Lx0EN5T8VtDv//rHC4RJWQH6epIM2Ti97FhiKaJ8E4
qZPFkV3TIvXlksahFjKIm7pG/B94KL1rEjqihWzOMrlLD2BIIgMZaTzcH45O41ONKNiQTlGa+d16
nhpHwMnWac+lT9PpLkJ4uRRa65bNAx5L5kq+IOew2gfD9IjnMYrrkSO05sWFx2nwpZoVbXq/1CJi
ydU97/nNLJC4GpfZfmjHmWTBWHJrrGhzIalByxHmQTyaglOcXE9nZ5Am9BWwb/G2O2lMwxMggZYj
2gHgXd2rFIl9kokQbUKfStX30D4CgbsuMYwzpHGSFQC89WOfT3fYUCM96+6nt6dmFp5NGsGSlPhG
I/QSIgWesKYqdogIX90mO28WJsO50/G2DtAxIr2UMFiJ4z8I9qReXdKQMdpj37VuoUb2yS19yZCG
740Lgdyz7VR60BN549hInzEe4ISpljCjwF7fRnX2U+tTmOt3axrtCZiIYpDz5qcwJWQf2yTBlBu8
32Zi6Knz2tqKsr/MoYi/GQUOrHt4ZP2g70bob7MRnMzbev0ekf4jSa1oBNZLP3d5E2U+2OUir7Oq
8TQJDuqydjxzql5zNcbKEaw+VltwAFF6oKIy18C8GBx3hGlocgkldj85qb+mAHAzzSwMQHD8pr4t
WS0V2C2f+kdztXF3B7nmgf8CorlIw4id9+I2ZHwudtvdiz/br++kLwZOGOMyscr6rEO1BoAtxgTr
qm13I3jMhy2M2mz/x6sHwRtMb7sH+ictfu2A4lOufSLSwxOG983pVe885zm0LszWvIxFapUO8wh3
W25YeKSG/R0Nd6K7FOSTpOx1CF2et3nPBVJmhpZC7Rz2WgGhCtcTF4jE6f3w+ea61Euif5GBwmPy
OBmfBY6vIEG6xwtgwgGYOg7P1QqLnLoG1FLUCmaMWQcgYhhNQfGseULUgUh+e+7iVq/ope5NSVoi
RRDB9Hw58U+B/gIoY7VwbgpuIYhz/Qmp35o/I1lI3vN8qVMYgJFAy7dckBMbLUEIFZu0d52Pv3lf
ql9NKEqjxWiUFWwkMiH8oxfO7GRipDzLSjg45KH6YadVbNiLYgyExURgfUfn63sVmxA1SPnX/qQf
mZWGcFrl3rqLEbKpcbp5UdVcwYJ6cogxMdel8/h0Q8vv0Q5UBHFgR5ccY8Upl2cFpppO8EFD5cKH
XiCXPzSwx+6xPdkHqhh3I4h+y9mBpoLHZ3a6zMl63RBj2a9v4KgyQ93xrMoPdyarS31NFUcfiSTM
sVwujNYmmkomll5LqPqs4e2eDF2ILN4twPHVXKt8gD7KgFunzWkpO8T5wZ6/GsMVOA0skHlynCDr
BqnWROD5rF13dsnJl9PZY+eFK6UdrH50TTiAlLP+9tbFDXtgf+t36KS3qJpjfMAWHNS09oagnI2j
EOJj9kZiEpNvngi5+9+fK0MNyr9oyjN81sSycwR1834awh+dfC5rfCa9vQblqkUXeJlRulCbVsIW
QOVY6XA/G7TDg502wmKtA0FNbpB+pyjUzmERva75FzlFVf68Jk1IVxl08YxVO9+O9rI6ATqHm7Fn
SAKQAsNjkBoEIFI5sP6qHyNRroaQUOBZjP2tuNqHpOiyZmhf6rYROMytMDVsZoIYzPRybmg67l4V
7j4J0FKM5k2KWAxj0MiwB6BJDcap5d5ITFp1SBaYUuftARefEeQ9p7HcNmGy4o7XzpmUw+RDtqN/
aUR99zxvJKOqJVy9AAh9G5N6cQAURfN5V/3EHHS2JQ6Y6bJfKTt+8H4aeCtPZypUp0kM9A1PXiM+
5uu4v9jeEmL523gWRymOHHQoKHbkfYSIuQm/sPDSwnBVj04lMydwlQZKDg5me6BJYufn74LNrKQ9
l/78ba7w53KtbF0ov6v5tLw++CCjLz6pvl1I1WcGTbBQHlEXN97CMXtEcsyvRDHw3UonvYdnnpu5
F6b1ONO7iV6SB2NMc7QF5YGMO3bLRmG9VjGMH8Z14SsUfhtcqKSisPYLxsQh2ewP1wuO9rFLYrqE
qkb4DIibO81mFczNCVhXfbUYPh0IMBWkvecSFOUjGJYpWY7wQopgPWcL4/yZXAzHQ5QfSmN5HHfD
79olIIdRDs2sozmnpjqs8Jl1T4nG90mFJfmcV4bBgXj7mWzzOgJxpPB+gcvCH5xEU5+Mo73D1UE9
+aTwEJb+gfseTvQHNrXz5oZF+u2pp0iJPg9gTpV3nK7pYBeigYFwUlpjdzD+SGiq4ihCDr/L8Gdp
fWHFMnCcwGGOtawLnX42c34UX9Rl3X3hEnT3GDGk4mbXInl8KWOmEcBMUaEULUsxxat/otJz7ZEH
rcUJKpIXwWF2732WWjj6FjOFJ3kGAU1b7t4PLYcsMfcFIsaoehXvq61Br/KGW3vFnhr3/G0rPk7M
ihFD/VXOyRc1u4O+ziuk+NEpH0wvf+C7SJncaFT5P+SS4oTirxxNOOhoIJMicTl4W4QmVcfOp+b+
shc/oz2JUm9610I8/54gSaobJ+VGRD3LGfKEFR8R9I5d9M9/cLto7w2D+vf6tDtrxIw4e+zzzBrD
8ILR45DLd7yNv2N/0aTKfcpjD1qjdhD1cjFlWbN2m9ei8kDn4x8ehcWw4EhkpRfvWBnpKKvUb2gN
NyEn+IwIV2u9AUk7xvcNEMg3mdwel1TP91wQl+Uu3rZYpRX61IRs0XOt5eErT1RfN8onirfFo46u
E2heugusrqxXYqDIa2sEKwPQERJlJ9qgJUkwPvzh//ocIFCStjbZGmRx05Kiusse6fXzoWNtimfo
LO27o3QVjtA/saTo2QhL2Hx0/VFOumkXdMTAVk6LaTjeCy/LBJvwP6QdMwqboKILhSFhY4ZYNfre
ZHiWAm2KoZKps6QFBxuPCTkJZ5dCYo2S5CMuT7Ukw0KYw2aarXvSO3e2OiuB5kfEe3K/L8PdxFc4
nt6qgU0AHcpRqNOW064nEgh32pzmrhJocV0PDSUsTF83LAqLnJKaU1sEJbzau1O/0Z9Ub7E90k6o
JMGqWltMjNMbdPjXwv8webz/gHjxJxM/zjGVKCq1TDlwmGPg0eX5KJVQTqVf1bA9Y4STEcfFm9fg
oqZ+C8i1vh3z5cp+lKq5S5iwkOZLXvOlmbP26Q5Za39PKSyhI8CT4/RWMLPtsBQCOT6XafaXIk08
UddOq6IlXWdljaU1jpYVFk3lODT31GpayicweuncS8IrtMvCqvWGH4qXGhPw10LSpS4/VHnKGtMP
o9hJc50yLErJa/xsG/kXPLEU4cmvbKeF1tgBS13oHYC5dgC+iidCEjntcqTnUBgQeU/naiv5BAta
KQ3nsr12nbVma4FhHatESryKafl+CIj5lHHR9LEsh2UcuLYBUvu7r4AKgK7IaEbVjolPB5oLf+Gt
TbAgI7Swh7UWtR5onJENafQLc/+qCEiWWfSFZyKXTjN3SZvxR2BrfsalFzzuzcZ3WhSnnCYMOH1A
VFxdVhDOPTSsDltYorE89nyAjt1TJKlXxx9ZjDtLqmM+5mfPuBoMwjojrm3q+sn4TD/4U1uU/BMb
ix5b/MOO+X5LDRwojMCgVqgFxu6fNTCcgD/deWtNmlHpE97FcFlVl/eo9aQHfSNn/+vjrbaVsk4h
1C+gj9SWbm8AichsrWsfhOSBPNhzn0iSKLeJW2FE9ht6VdeklM0aSjLoE3WTS9H6RjGqnzvDntYt
pyIr+kT0s7PGKADIpwpiRaXAE/dPAjkkwJ6+OyAtIoHIlvx+OzhB0CA7U8U+O/mNyWfNE20nmOrp
SxwKRvv1Dy3aFnjhTp6SqfiR7nRVQmbcjZx481dkijh8iNCtBAr9R0Ci19lhufEj9mNGd8C9VINv
ZGruSJXJSeKtVU3MZ7sgW92ThCpB5CIlsHl9Bij7Kcw1HOfINvSnzCqF0AiSS/0eaW3CoP7ZL5Y2
qQfiAFDGW63ECHQam73lWfK2wcVF7QyoK71C1A0DJJAWpHwBD8bEGXUdO39krDWWOOIWIwOct1di
tcDcSGFkInwx9fzDViMlRl+q/0egycHEVF5Wu5idlzNS5Eef/0hoiaZnUTcWcyldLNKCFMU8Ej0P
01Rxw0Pvks4UC1aIAMEar/3yEr1U9UDTe9mYIc6Ym0KeXe+M4xFj4XYehztsZZck9pbX0lDJebx6
jtw3exVkl3J0VTAO0sx+9Hqly2B7KnkI0CEvXfRkeW4hA1frQvQZj4kzLNO7d0FTfRzrCkBjFv9z
P4hc60flbQIPPxgAP6mwx25lb0pNCrlfvtaSkxndSMYwxIg/Mh+6n1Y/rNaSlhQrXg8bk+NuhyE4
gFQR/e+/Be10uqX43SAPgBDc7C8YsWNtCl06AIhjxDNtgdek1GwS5mfq2O2/uOT0oylyqz736EOf
bytkqIEF/HhgqUH0coiGxhBua/ZlC+spEDyP2QrOS1hI0YOK0wTsFYr5xIH2p8OvO9bfoaeMwiPV
gACqpoN/t9aMNr3AEP3rWiVnWTw8iDUonGa72/Azdzyt+ejwoAkC+IWulQ2F6+9miMI2og788+iN
yMK7W0EtWQ/A1ukQwU5ApBIxh7bbj7qcrsyJAAmpg6nwec0tyCpBRTqYgWykBSk1LwlUo+6LNpKZ
HGUs7UDpktrTxD4oPq5kJ1y2gT5Xq6vhetYNDECJytQ0isTLdlausNSN4GM8+b9MCLyLRWPkbnKh
+MOrUCP0qLu7jsy6ye5cqs1YDrpu3VgqIVNRhzjP+hU/dcpGumQlMjF80Dh0EWHFvakrNF8niNgl
ZmVYdYU7HvmW7X6MkCjwvylV1yOqO+QHwcOivOO4QDSv9m+NSwq989J0o7n1eGxB7PhQDE/QSte5
s9W/bZvoypY5n592mJmTA+K83+UfKErjAT4U3A2+JiIkzfIMnAEeySOmalScxjSvEiVXxr/ahMaY
qv0gagvsl/GUIWBQ6PtDAaLH0YuGgDTLwswCPoZ8ZAj7/mE9Ny2yu2W2qq75lK4AZwQ/TyZE64+C
pln3rrPfNn8OjhVMEkc7Ab6SAC+urNDVR6PAlAg+Z9sQMV8aqZo17OKOPoJQPF2MmA1ntO0sSXv+
PorZz663aIOPCmyUiCPCg7020I72dLfT+tvZga+RflqHL9bi2L4OGjkX8e7MbI+xyACrxxmiVcee
5FvwN24VC9a+6CURiuKyL0WnICtS6W2BRr2Zsh5cLbPviVwZEriGL2IvEwGm570ROvT/DjUVLj4f
iS7hNpwCdt50s+M13VHy2EkegRBQGBXp1yjpEUphBATvxgHIYprCf3DHnErFK8+Z0UOmVTxeacEo
s67TQvH/ePxtHO4jDfUbkbhnINGi6pefV3LZ9EdxJrALVvhBPSuMl5yUtaZI3WCs3SBUaFFRZNyF
lJrFH3huSCVAD5RhxQszVCIzEdMg5/xcdglWDwEdZBwi6KvXUy8O2RfRqdIfCFZXZQbODVZmsnYM
ws43XWJDq6PFZrurVdICLmehOaI770CA1J7JJn+EMZ/VG2UEF7vCtujmSDgNRiN8praD2RrsMSNB
K4SRw4/01ci6nTFFyoCWD3PLhBwS3g1pKscY1hEe+2AyYZNrMzHWS2UtLkd1x38JWlkdLjBen3Jg
LPOU6gIfoaVSgUSgVqrPkAr8MFn+T3tmXm9P10Ekt1uD4sqDZu8hWl/54RmZUMA2RNpGn2DVSb77
nSm21zUmavjSsWv1cR6/gVSh0oh9C8yh3mGUdaVT7eMzWTkg8q9voXFdGpBYpM7kK1GjNkUQVia9
GbgqQ4P6prfEnk1l0x2CKe01q72A7MRUyNTi0+bq25R3DdJ1JmZM9idb90qIQAgz3pPYX2X9Pjoz
AEkLfAhCYkv6vR+vDLttMu0Jj7j26VeCSYl+3ewUm/WXdf4lCLMYrU0eiCQv21pdW2d1ptn+yNiS
uR8o5ujUMqhcHwwwEYg7gWQGVhDZGbOP2FsiNW2SedWmI6nZNQ9MWL5aifnXVi3/xXTjMB0U36EB
R+cZyppOddXEJsBBcGdorNcHs4ausbr0LyUX63SvJ+LuMXy5794GhOvzzZhqKG3g46nE5jqzJtRi
IGjA+qXHcDr4BBMQtr065/9vsjIyD0UrpNIRgAVnPMlUEDNXEyboFW5elC2CdG8oZvQaG6Cgh5cd
zb5SiUea3zqe8iA299Bht9j1yTUm9px6skvUxpMHm5sqILx6ySJeBCmfHxzepcY/yucx6mc9Qp5U
FsSL9bZDqkLLK9PExn4asHZYjiueQXyYciyEz76a9czFo0q4W7K8xU6cTzOIXXoh7xR5ljL+incV
A9f+gEsKdalrvd0T/hzS0Ythk0QsKnVjFb/+MG3/1cyeexXvtvWGeYewIHpi64VmrLpfAD8gYPFB
jTNOySITdhuhJAdRBJ0aNmoOS+bZQYZRs7i2byBa/nRJMaUoVrQhoeWQCTckmWco2JSqd9YxXQQL
J5IiHSa0D8l2GzvdMoSmHSZttnUSKL/AHSeVGWocGErriHt+qvxNyze56G8aym9uFf+AQXUt9Epn
lSENn5YSbsiMeJIhJFkszvwrn7LNYu72s3noXSyneEnI6n4e1bCFfcOgNhoJXPwjw3AGFcqiOrAs
2U3I+grQBGbqAsMRDFzpp9RK3Bxd6PDlk3XhD7RfvwTB3u6A7QyCm+7xUIX/yDzqeCNRWst6UqRg
f4WoKUlLTQrQulFD1zHcX8urSU1bPrj/XiyitishTc5XvjIi0jWzQDe2asaGf42+G2tCPbbqw7cN
FiYI1VALJ7yInBPJYWGq+GoD6a5j8/YbgmeXshgWjC6dfCHQXNjoBRfU5SbSHv8KOJAvTUY/wHUt
Acgx/Ic0ZZOLdRElg8A70itCDUI/azCx94Q8uOp8wba/FAcjYteUxY3TGtqxV6tSkSo8n1n8d6ld
VUXAdC8naW3FnAceEqm20MFQSoNj7oLZ1nu4ZCuY9FAd2eqns3H/3d3wwFz5SJDKBECRFoICGsy2
MneiTf1V/xEGrD1Cl/GYkh2PyHeLaQ7I8N9iTkNF2V0rpSNN/2qiB2bkIJ+F/sFq6NV9YcPkYswH
2pmjor5ErtWSwWkZT8bv3GzoQF2LCNH7eL53A5M3Q1wxBNPA3fqZBEQ6z3uZ0yxPrTOtnJD5/QiL
46e0Chg7SgJI2b5F+aTNhITK0TTZmR8rBCj/CmNTMVkBMSp3910/fBAEtyPF/7o09XPWKjDLI9SL
DDHo0UzXwQqAdEZXubAqtlVl7w1VJK2Eko9Qf3XMA67BkrL0LAhC6DFiULEKLau1hhYffOij2mXT
vtAp/P1KL1FqHBfYuv0oue1stFm/5uKHvIM5tOGJm37bHMlsKcqQIcwTp8efDf6SdvTs53uij+eC
yiGeqQ8jsxwpNPIwAhQtuY0daos/O3+rFz8lc67cQvXAZLuAJcR+dEXEjqDkcPYj+cRT7QamGwCN
BAMY8bcCttfmcqXDflZIN0amBw/+V1av6+1g4Ji+PdqIFOoYXQ9DPyaDTNneBp4u2FacRVp3WhdE
jZt2Ve1LzQt7Awad/cyvH4YRMqanRu3yyBzgUS3FuAs2H1Hoc9wqcCw2wZ/bveb3gQgZUpYv0kZp
ltkUJfDWjsoi4wwFTJIM42LSc5cXextaxIgAcpXpR9q68IoMlunfp/7+6403K+mqVFriETVQP9aX
gogv4KMf6PVFbzOIr7fBS/pyWzbcumcVdNdT+YKCgnBuYEnzhhs1udd8crE1Q1yAPQQQ+0Bw8gxl
N8ZHCpbQdJwmr5+Vk+ZIAIAQLI7bDiC+YhqGZojuS3QFusRWwQ4FYelfcH0tu4X2g+bf0k66pxQ9
yAVMhx78mElgszwzi0SEDoiX98LTSPcb0OvmK7puR/VDI75AFcDB426+GGgp33oR5P7Hjm5v8Pjv
a5aupPSJVfXExI/00/+uXJ1W7t9MvBmIbxxObRwfu643Ta4pSlx67XvJX1q/WkICz7OKOCdYbXQs
s2rUcl2eQ9DdvzaTGyWdjwS56NUhJEgCAwFRjymMvnZsWEMqljkrMpoMD7kxZb8QRDOZ9J6ezuR2
6idS0xmaIWGwW3kljm4KxMVvkofvjIIpiLcGu35tuKco8Ejy+o475MeR2OllmPuYcnS0Fy0+kLYV
87XdOTIj3+PhHgXlSllHQ1W6Szpa6bgHwEc0/yt6FnQ41yjAOfOgODF77Oq14oVYhvZHYSVWtJuT
dTp1fdJlAzsCJ8NNSmTQcYvW2H2/IQid4JMNCCZUcHROsN2osB5xKsVKI3GAJLqhoWSApkADRIHi
nkTwBtBEIeZnztq8hDx/OMlKb0IqCldAbiR54ZtOLHgpJTF5jEnH+3zMYOUB9/z3ESyi9GwTQGUo
HOUy94Fw9fdosuriVlTRtjhw0NIUoEnT7Q3JO8IunNaes+jEghLePM87xSUWnDwZDNWtBupixNOr
XT+vgFZLbPAj5jAuSq9wPydSF6j8rADexexPQgLXFjFCD3eewO/WuDl/GBkcFLKE++THtLER1owW
Zw3PhaKAzHpBeDGb+ORbqOLelb9nshKlNF6JAAkctkAYobmfKNIgmnt+j5/0q9k/Qj7+SaL79XO5
2tUEA2EXAV6kV7EWwBEM0OFhcE3MxbuXmXpOMKNlERzMyGzyCJpS6gzJ1dTRvfBwkL5DA6jjBhqJ
ZlzbFT3Ybh5n4DoNwB+vjNWYWYerokmQ55OT6rh7r09L7UeQuZ3/k4JHw/BzoK4gVg6FiQf6Z3k0
wg0Ni7iMTEZNs730slkEM2VO04WEx3X7nczmnOWa1CYX+xYUr81GHoAgzGQqj0ejMR1mWvD4NOZN
0qtfql45UwCMLEY6Oyan3RE96cj6uirPlyakER/nrvEtPg38cEpBp/02oSoPPNmj+NHJOiDB1Gy7
SnJzMnN2zkfBW0JkIeFDVEUzkOy3TVzhlseWgvnc/GiNiQHyJsUjpChF4fpymTf6bb4mJH2M0Wrw
fsPpnverdjQ7pz3X+UKvkuAkUtBd/7L+QapAS0rKs/TfgVJmvzrZtymbiPQtjXZTsWTaVsolXTmz
FqDriaax+NEAS+vNrrRvvmq8frLK+8QJNR+3KL+aQPje9aDzB5PJy0TLBS9hv2eBI5YIOJ1wJfeK
lfjFg7wzaCt83PTvKX2mQ7BwgPNYuPWXBEL3SDCke/nGqZzkveRcBaQvwy7Nr9P75Kq339wqEmLg
NAi2s+aurgoU37z2khAZ7KY3im9nGwbVgvNYnZjbKxm62pPsShkDDEkj7v4eJeAIuxd1+EPyTZCy
xjBkmPIMy5FnKr2C6gtfwurcpRTrKlPtDQSLN12AC2TwroSjRZ7wjoSFHGzd6qYjC5nv9PMRuW0u
TwfGfpRgJ77ouHruC8p2bYQuickHAe0fdYLGJwBBBlsuLEQFUip52Yv8Zgig6ktKnV95A4voEp5s
o9AWIV5s3retK2Q097gB9rLWZ1YHFiHknM2G8tdRggHyxXRb9/EEUckv0NQHO5rvodDlPRvMm+aG
BFHpDNB+kP3cVd5N09rVzmMdFgeNnv/0s0j8sp5otSLJUosAWZWgG/J14TGFgejkXvqvkV8XkWOc
EsaLnZxsGo54eOCenGd/KyPwJKwANJr1Wwva1aGhII3YIB4yE96SoPqCJOa1Cd+mrHiTELX/Gslc
OedMd9QYO+x6KNzFrqhyMUgf3Fw7oXMiDt7K7bBdMawMDtqgTw2cuOU7F2oRncE/rnuiB3YLdtTd
IiWZCPOew0R72y8exoXtWhI5MCQ4rf44Im/qInnuWSyb5FHXatBd/FtMj+PLj4RinKJxTjCRXBqU
CsTdonHln6sNekqolscgAwxq9cPpYbVg0M9cxf9Tr2h/jZ6ZEAn0ipqAIVszGQPWsZ5NaOl7kDL/
OalcJp9AiWy9BoMcLOvLC9x1+Zw7tP56yJtlXAwXx1VI9PEJayMUUfptzGGJSVEFq7W1SgmC4WJ7
7ZKXbAP9bosnbLPm7XiBirRQcTnliMonyhUYi7umwe0dbEEjoXKPNKiocquSYZogQXnlYxznN4ba
KrBjmYgT+ugXT0/mkdyORew5UDSP+K43k9YBtMoGJCNBae6duCaicqUvc5qIjtrsy8sGKYqCprnS
FUbfacXiEbNOLNkQ3y3Ga3isu9vcdgkIrJ80jxLB21BCPpIdhh29VacK8n6eugh1muQGWac2Kpzb
TCzlTGDqOqoWVbCWEIPC9Yd3jwze7/jZElueGw2ovC9iltODGdkdxuDw4dsn0rs9rr4vw0cAnsTV
L5Y7RLXxAPzvOHUIhKKx6d7gmIr6MUvrLoSjs9+Q6XRuQsExJmrAO/5NAQhvJchmwdURn0QCP05C
FAQA3q3zYP0Uw8Vgoh70Ii0dmqimbLqhcgJK3PyzGHKAVMbKzweknCNGSX/5XY6/MJ/DGfipxkZD
QH3WM4B0ufohwLCJfnjynkqDIB+iEDAQLmzGz9Z+cwJOKPB5Z9Hb4FIYcLXDaSPbMVxNfxPtjGZw
XSCHlArlq2F/2S268jesU5TPzlSd6fhRXhW7ihIk65qv/ih11XH3S917+QLJgB1BIR3FQf2f9dyW
SWApoG0poDeNgA82x+lO8t6/xC/T3XNP6Vmwt3xVUaGhhZ5E/d4+XCTyQja851lzmXTN7sdTebLt
fTirwYfI+IQEARvZwSLf4u1uI5qb9i6Qp/jA3y9SQzGuvaVN/CuaLniXndHOX9aHFD3CBHo/XD7S
Oquh7gXeTXKEmVmGe9Wr0dRp+dZljJUa2joxlJ18gQLUo4ZSmew98tD8kLAM1vteBWvt0cBANYSI
cRYkVnbbR5oHylVAhGxFPzORfeydlQ4H7vi6GANsemxm8BUtG+RZNCl5hkG7bsKO9R52ibmdHtDQ
Wila8Av/t/S9wMk5MNJB6eW4sXqBBCbD8W0Sb8FrAbpWDhlSM6EFoxQGHeLCogcGkbhVEk9/LRYr
H3SypDl+BufMcM2jJftEybozbQMk/sGFVHAyPqe/1s8cCwhWmntfrXnGtf3Toy6lNbnIsU+TyIxo
zW0FjfscQs1say+VrZ6K2MkqhQLkHoHJTXwrmOCgyR+0h37L9X9PF+cioCHoPH/kMx4tucinxoko
Avc9GD2R9wFYToew+1UbyCXk27Fa3ea5VokT3IQ7OcyrwdSMPOxVjgyDtazuFZj8vIgyqEIuRIjw
okPuVyD0vPIbI4k8EmH1OtYwU82rZ3x18lfcz4il6isLeivSdJCe7Uz7KwcRxK9caboF7WbjZB3i
xb86yQ2IdTsbfy7q6c2plT5hOZb4SKq3JUqegIfDhVXVpjCGDJZu+hHm3bidkqt7Jxqbww6uC67q
/u3CYTGQTbxIzcSCY8DPChRspud8djshhppWk4TD8aiQ/aoHH7Biy57xPLscocwUdEvlnp5CGEj4
HX4rnQ3JULXDXDS6hTYbAL+1+agTaN5XtiZtdfDDJ5j/Qa7x9iMBrtnEj2Yl6bIeuKlaVnDa5adY
C0YGDubamuglAoUYjh2XKG67cCUHijctdkSvKOmPZUIAPX46AHDWyARFwZ1SWALKCvXMM9kYHdwE
IMyEOPAvwLlnpLvOk5XWvTPxXnExU8T8mTIuucBXqhp6gMLLk5ZeFyliWM+HCTCgp/aJruvVbciU
gNq1oPvIfjGsTt9lDS5x3qdbu8eRQE8ID41LCb/MjEEGuuaER7ekF8SJ+9ziQ5tnhLNPxugdbkBA
keq7lHCe19wzgdmiCQ1CCc1o5epDNRsy9I+D++og1s6lwUyha7NiDR6s+vjBE9JGHsVKthupqxXQ
4y4//f833UQu3ravZ5JL2Vm8fmUDjZg+1/5zhdUHrd3CB1kNf+1TkuxaqRTqAGxIxx1qlVHC7ffN
KJ1X32xrT2B8x9OzD++x4cZkjHIaV3hcQEzAJNkyOBDMHNLJwE5fnS47zs4huJcvCs3oElJeQIP6
JnOmFnOi31i/bSit7dwRaGZ8EZeQCkCV2T6U2vbQWX+VdkiB6xjgJxit8WKnVFFnHedETQ7svabK
Ju8TLe7mnZ4nWwmfDJi+Y67BLtPu69jvYf9wyZc7UVhR6PWkVrQvZU9WsKEix9hSP9GpdGMLpI8i
KRb4GZ8k5QRSAetp3GMtBO444yRhiYCUyGKd8W97xfXbs/QuhK9sfZYdpCnfLwt1qpYm3rjOc2+7
P08wbJ/WetBbCGCQ5K3fve2eLw8LhLwaD3ZC9eHUrCzkaTPTsNGR7+mevDZbrZN9c9h4Sj0cGUGq
Z5gg2Jo6DLM7v/5eehua9vLjDstcayYM7emAu+H/UmbFgtnPoLNHI+zZh1bN2mEKwUyliHjRjVil
4lVSeseMZlzJMaihJ0K1mqmfHVT8um4CapbdWMzdhg2XiDrzqpBrD019rZcVqSnR7y3Mb9qVfXgg
7T7N/sTA37mKi4knpRb0b/mf7N9+YvPxfKjehQFcNaTHwimHSs5I3BKhi1g6LXeItt4gadpV0T+T
dJ3ZfYuTpPFkZGAJSm7rR1B2lLKbYKQ1axZ+BqlI56hIiw/PIuMSIGWt1sSzqfJiQaxlavHRHIV6
5BhQX9GSiVJU4AfX4457Gl/2dTJzvKNwBproldWDiA7CtaqR+s0UFuEeWAIC6NvClpBodELVuxyj
/5Sv5Yj6vc5bxtA2NL7oQb8LOuZD/yVBF2uTYNvma0MYwaSD4bpcocOZ/GkqxNkwzmKaaMjLjzF2
U6ww2gyjUIYTHN6ak+/mssB5kXjIH1gqoAUxGbtuoq8EyE8zN+gGK9zPy+6G9qyTWp6cm1s+UDgr
C6BXiOKYEBdGB6XtwL+bPujct83eSiM02J9932/5VDz/COiUSagkZrx+zsipnl5a/e4dHVMtluqC
jEQcEtXjJZ/8oykHj/9ToOUlaDT2FihTkuTI1L1yZeyoEeedDcz9WJH5T3D3Qa4VQrWO3QRHumc5
qyP3jMAeVsqowyyrsQVE40tmttnJo2POi9P3rOad+In5QS//38qviX7UTU+CXmEVDG8N99IDYS1E
IzikuuP3R7U0PKUzXRCwyUpil38fowOC4TSlZ8rsvl7kcjVvNm08aEuJWf//172T1XC9qtVIlmSu
6WlYpKzfARM3fboDesEloYrFq3fG9bJmkO9FrIcXt++/5hUbpH+k0xgtk3Nzpf4grUHCy5M8DXmI
z1BKJZ8eM6yfa7KTckaXAMqThZI+z2PslSlbtObO8YppgfRkLIY3T5Hkv6lXBSzbrmr7TClhPnI4
Wd7nbPrJJDr/qrqJnaJ6sCqneb8CnPscVx/u0r+/Fr8lLqFEbsKkAuCP5gVGTsEKrHpIiSyuj+Ol
+SmhTaoufilS1Bb/OfuF4stNbk8n+ZflQ2172WlX9/hHIu28pAR+0+rrfdSziJW3K7p2tmvnRnHD
2vT02weHZSvsLo4Kaq2sCj+P3RFJFKj8PT6c33uZgzoINp6ha1okORrRKa911BNN3UfbfkvwCt/5
/1pryWWdEoqKJI7qfOGjAjKo53If99nj7d+BXIh83zJYj3S0rqr5jf0iE/EcfyZKdbkPNEgbuscp
0L4y0kuKq+GwmNtpuX2vZVrYkkjQqhqvVtR/2T4pIKkqn7m6KFvgQEyl4uuppmvgzDQU5fn7A+iN
/KCF5mC+JMEn/4WGKNUoQ6hdno/0Il/zOQRX73z/snaXPTsPCBik1gWXKvTBxNl2JEwcmPGE4fNQ
Sqard+4TLrDleXWktAHT0brW7gWn4JJREayRxbN2vpbrelhn4pJb9MLPcgCLhjAQFI3Ok37lPHzh
UE9MQhz7PGIVx2qeQVLV3dDkvEF3NsxtfnU0/v2E+j4pHbKvP7ZtKzUYJzCRP2+rG9rW7ILBPSKV
8e1QGQl/xsXKztkvjCV83GC8T2dvWj6xBdCUx/j1prgmtyx0tkGChsqzHk2gJ2PCzUtj2GH7fj6Z
Vwpmvqy0rcX7OCypMaF0rHUlEhb5m6MUezdVYkUoJU7Bk1vet6trJVYExMiGuvEAAc/L3QaF3amm
1izJFEvI3sC9pSWnS7r4Z9rQWmOllbfyHlnZ3HhZX0bSHJwW5Uny9I34nrkm50B0w3JCfBsoC7y2
1IlU3pjGN7MfC2D6gpeLCEJxEIw7+AEDEZqsgeqYX5HTZCP8xbeeDrnRSwm0ikae/MIsastJPQgL
rLst4uU0XrB7XLi837n/dik7AmUUggl+4vCUubn/F/bNiuaiXPtKB0NJ3Z51VucZZWPuMP9KMVWj
Qkd5DNvTHvC+CGMeEazIjlBhdp/JY1AtM0Le+ygxMkzd6wrPdK7y1NZ+GmI64bcT/jN+rg5niNzd
IgUtgIr+MepCaOwTg2kh4YbO0Vu+ci4xCeArOy8di9zwbtq+DhEaYGVMI7x3Y4QHpOmi6H2yfUTL
frKzpj2hWtoXAPxCOopIDSqVyutSMrX34TRJdy0ZYTz+aBtW2686S2JglzhaYCdUcjv2YIraGYZB
mpVKUOfEj7alZ0uX209u49Nl1NBGqUozWvcjR4JI7QyNqcWKG4ZNf1MUJCC1N/bu5q1yT9MOm7cQ
IbHzae+azzGZ4dGKZ6G15Ci15iKTs5MFw2oYJUnogn4I8w8GIk9Sn/3aXyMBr8z3xkK3Au1p+WsO
CeStgD2UbP0UkINnvtr3IIXUyqJEsPRc3R8va+q+mJcBBvjgkKDw1PFRPvG7sfHEyh7yJ8GHJQSl
OrOkpb4vA0PBLQhzyDrzfWRcbJkImquZRs/iHcud+Z1l6DIYF6USqPTQY6UaXm4vplmZciyCXnLr
UfM6v5745AZ8N2DiDjl9RN3Hf3LoSG33HbU7PaOmElIsw2+5bjdqjQWtEbh2NXLvuHNoCspgbblV
BIGhUVDgpMPfn2YZOkWLGQhQvAYoHMJDHomxpjpgtBH/tCyRHbsDld742sFqe5DnOvWpE7cu4SAb
BtfFFnDdbQ+kCaGnCdU+xtrsxzLUnPzgRmxPpb0PlwRLaO712R3NVGP7JjzRlz6tHmBKMPkWnFvH
g6sx0dK4LBn1vjJb2MF41tyDgShJudpmXvrEFPHgC/XNOHTNfw9yD/AXQR+mEQ278qdR0xVU2wPY
Aw/8zCLZmhJw4bL8qrxsYaYqJp83DQp6aAlJrFd+Ted6Ny+USdvHLxUuj81s0/7ozSkoVMHNH/91
CVmax0pziuHQLjsF6LGKTK3ANVqZ3cZ8X/wMS+v7FCxqFCVlHlfynxIuTj8ApvA+9orNrAnxOXQc
4hERLfAYLvZSy0ciIQX3bcaO8fUUzoHIoDKNgWvH5nNb4OokPePoc1aivC6H43G58ShN4mVjgmkZ
CUqmsJ/Lkn9ywhNT2zzlF3PQ0ZKh/GTZk+6l02pVG9u/6jGVCMQOIyOLBSorWoRHwCNY/YnAU/sW
HaG/Grt06pg4f7bv2EcRcr8ZUlwLV5/ttRFf0pOalEoH1u8mQELA2L+b78FwdBOxrYgt2hUu4Nfm
HZxjLseoRbQAH/ntyDGaGuyGEIHroZ9rXKgYQgxUuaihCDKwcAQe/3vUXu5xxXYGyvw/qY92qNLP
okNXkOytAszNn1bamASZprUqASL0K1/vjyB/TkEmPCMVr2dLGYaay8BOCsatZCGUSI02ABJNB5eM
aQvx6tllx7L9k8TC3ITPRnoPTWhCHe6ktAmU2Df67gzrH8DsKeuxYNsHNohwjTYtK/I4hVh+QP+x
DY1nuHAOGt1/16Lq0FJbmG/Lj+ptIV3qPkwh7DU7dKIXltfhd2s2gjalaIUH37IDTF5pingUKQ2e
AdiRkM3kLK/ewRR1Bq1TbMVFedweoOsIXhry+cYsXnYDrN2rX7fJmcw7CHAE9j2fLniyp10vS9/U
crNfPCgSHaF9CiSSLU/uo6h6FfWY9cIzvwdDpZcdbCvhuwrprM/OSo1gd3vlF7uVCJ3oF7ztv9X3
wunGapAp5VaZc+RqHKTVVEC0aP4pMN0aJWWXjec/awbWIEN/IF02d4wl4DrZGvxLUTZeJ+0I9DtJ
5uvcjv91vH5Qyp8m0aJSvp2y2JIl6GvEkoqj277dKDkDAkQoIhkYrfJiwkQBosnbHdgYpB2f7PFf
A9uGxy89DIjAJpmWYRt0dnJ4ePNo5nYkFz/T55ujUVYfkTLuJfYcqqQxicZ9e1cgA2DNrmYobqAx
QCZk0i0dj6KyNwYqooAooBzTv0KEJF439zaaxUJNYJoCxYtc5PhgIkGhyp6kdc2S0sbcjYPKW/Og
I02TZOXM4iz0NeFDGvjh30PsX0X1yO6VJrZaPBuW9scTcmgNHX6pmsRURudadb5gvS1gfeFab/Lq
TOL1U/X6n3mu6nodSbSkJymxD08Vd4OMkvK19BhS0tOWzM3sYbXAERvRlCsTvb05pCD2cx1dL6Ya
whbhMBLAnkd+QqG0Gsy2IIiAIlj5cwhNjQzFMR0gMPl6Dxik8bcO2lEN9N9zqQfkZZSDaDqnd6Xa
LmPMzY5P9KIMWi0AuTwvTbFd/0yzSxk7vzf7ZxQzXtFF1WJgdji+V/5n+ObRT4BpMhzVjt2g2gM2
p1QgEl6LjpxTtr3bhCT0Ah9aJhhVcBF339L3hXRv26s9hbwJBMQrbBi6FT0GQTITlJYcc+iMBBcf
W8DAwOOYWRscMG3/D/C2860Phwjux76qrV0lV7gaa/c1RjEBRsaNPW7VwxYl6Gsm7w8wMuBFqTTt
kucdYa2GTZrA+WZvKuXuQhwRncYS83FYlguvtP2VxTzNPtAvvE2N47IQ9gpglhzTg1LJquU8x8MN
omiXsCzJFG2QZ7o3o7VyasTKWittTaUmAj24Qd9NwXySW9gsHW0HtrqwnNjVn0xdzp+EhGE0Uelx
ZlD9fC+jJvDkn4wLhyjeTfT/YJWBgMey+El+6nMKKz8aXjtS80MhD+11uJBGbN+A+qIeE7CBdN7A
5Uu03waDKZ9y5Ev1zZToQdOEpEDTKeEeujbIrY3sjmo5IGwiondqzciUslUl/c6wPdQXVkCqDSgC
aCDC5AItgeeeIeWGgbEPHV8REp5UMLDQvA6HaMCpn/6PuM7wUkbDbNk/cqjqoOeuJc8UEB9kO5PZ
R1Hqqjk+5MSyd4nde0WN8CA3pEvDJoHUcWqNTmx2FvtLVltdDpBzzlnISR4nsIHd0zvFH6037pY7
J3Kn6jMmWtmVjUfyfgbPs4TJVX/qGwqCd53s0gSdUEWhgHtHfOfY08t8g0P1LD/sYsdsgRTinf4C
pqg5Wjfajhq6NaImXHL8LLp7d13LkY2z0tqHEWII8uPs95I3dmkQILZKsg4s5t4Sh9eDN+82fP0g
x9qv5/XXGLsnQi86ZTt0gCotZZozpgSrSjgGBKFC++4NR77jztXrGzGK9jv2ZjFTASZLKe9jp1hO
vN7Vw+4e/9GP6wh7d9XLL8I52fyPZyRmoHEML9QoHLHLuCqC3iknLaMwAsG5tgOxFY4wYNsqDY15
aPiL0imYK3i+McxnWD5nnHuyCs6SSM2BzlpbcvbiFjubWPMFet3uoCHzgGOnFHZQrEaGmpfMblV6
PYjQhxU4oIntXGNndfG5i+QA0UXb7tP9fGUDyUQsgfbD+cWpY6vHF/p7m5kFo9QV/XugSl9iuCrH
OZYcfqLujevTTQjrLZ1f50ckaUincoZnvR0d0NchoMxwMe+D9fO+wYr7PwBPNVlDDBMOpOSCwbtL
amIBf/6cZ3VSewc/GUIPyL94F7t0NS+oLmb+HJt53y+fgZA2GVjCcXlhNVUdjazuK8kWSvz57p0E
GpNpJ8NFi1y5KEM8rsaZAjUt1XtB1eItrr9hsSSiGVjUiTMIRcd9DfMjheeAwMiXo7auAnyfKkbq
6qDqB5MqQbmAOIthBo1ykdq47Sj6fPr1wTZXLy6IJ694ZR55LW8r+o9dKTxUAi7354jw2rEF/NIw
GKMYkV20guEBRFqX2cPoxaHZ0FdtbDL+W9H1tEwHIZJyOrZQturraXc1Sb3g39l3ObJO3diVivtF
K62OGpRBCYD+8vG1elbzAQnWCeVUof72TFuY2BINdMvcbZfaxKhe3DCIH/YKeTZAIic8RSYkrzOr
kZ/EQvj/KvVg3NEcP1Nt5MIMzcFiz8zTkDffOQrZ8Lt5MgDltN5EZFgbL5Kd37Q2IrQqiqgW2iug
R6nIivfLjL/B6JQmWOK3im/EDbgfb116E6ALIVe3DLVqeurqkfjR503KnpzgdKh/H3hGolWrOgu5
5MXB4p19HNi8UvtK6l4mZkoj6zzggO7FpHcPWUQrxrr9hOzUk/HBJBkIIRgL/D9Y9fKNoHjlphyj
KC8d3liHnESMJ1OiOvoM4A+nQFLaTVYq7YgXaLE1mVvEIgfAp6TK7Rbd9buihtyx+dz2MHpQx0Lf
/qTCReaFeUpXVR4Wb3MUw8TCOqt7wLNEPk27Hz13qv4uAPAiVIvDptchR1IKNi2SDgIIuLgViAlp
S4/DIJEctYGHfvgfPpJ6ZtY5g6CgxZFuZILxBr0vf63RC3AQ9rqDCCbs7juMzaoM2deFOePc2KAR
nByAmbal8DSP4XwoKkQepTDo1OBDsK/qGDEFBX2Cw5CMFodTeoDmEtGjQqS4dMewa/1tc9X18AVR
mOBh/blxQUOjH1UDe48qJw/Fvdqxs4pPlWScBuk3Apn9xp5ex1cQS9fIdIQXwYW28wC9fujZaVLJ
Ej0VpQ0003OEeaYXAEPT37nAnNzFbjdieEs8zgTBNfP1PaOi4AbL1YYvTr2cxIA2CHrXe/8SAkFs
44RYI5G5DvnMpPA0TN6yTx+/p4qqGwtIMXpxIgUvQaCBeZCtdh4E0kw1Mev6aSqXJxqbrOLgpc2X
IYXCcpOM5ZUPgY/Ipdo6T6DaaINM5AKDaIaCxrfk8jJgk85GG6Rjf6q+SJM4lnR6QJExdFssvETO
MR9sIp8A4t9jZqJhwB7Yvsc1vamzAL4kw1EDipHifHcUieUeYLjUxJpPJF2bGorFlKZ2y/N7ikcb
11GTOkRlR5/vKGA1xik/uWOOZll+l2kTAtFFhCFtcr3z2Nn009Nj/SXvY5jvnhrtlZU4Tia4YukN
N1SJH4PQolL3RNe14syQNAgquklT1r64L4kg1yi6DUyDmCsLb4zNOtyGuABJgUcvlYabHIgsRH2v
4bGp8SRij4ssILRoV5f0NdjbMCUV/rQQzvGMAsX48oz4XYTHJL/GV8PqjmSMUKtseInk8FIjkfsB
UM/M2WtFp3W91PhRGVeHgiD6aB7NRFQvhZsY9nS6GKIZjusmy+OH9krTFpZ2ix2qs+tghrSWV8DP
u17pRSWQLxAdAgHDdKgYAJi3w5uUdiUpu8MV2QKhiV2lREEhsBpqb1rj5MO5oqSq69sDfYA92HjP
XDGqSUi96Mwsaara9J2D9x6RA2sebPIy218tLWtrBzFwKf8EjODrAENO0i4X5pbxeKvm1oOYQOgS
DsCOkBz44kULEhvp07aoHMxRme4Gn76aBk0snhAzfCy6PWyjSQsaaLlxp817aUWsabxiaThDd0y6
ZVKWp1ouTRXOOJMMgQ7cQnJTlpKFJMzaiSGbVjijNDF+dEQRFt8dA4gTEUqtfUCakGnEz6l442T+
4dY5mFVroOMxIXNeGJJBXCGzvgJWGD1kW9sH9RxTT8jWfnsyDa7RNik2K7/F5KheO5j7c7uQ2Pnw
51qvRyShuuDSSbAg5nBzeyHKoUw8gzA1AedO1o8psyDkF2M1fddKoBA343UfHSZIfED7m0LHIDGg
NbGqxqjEvwKQgSWevTZHPQvViebKx3MCYX9knM1p8POH5lZ+3BFr5t9oRUmDFv+DQ5e80kOes3WS
BzKlyFAYICmA12rwVphdQSITtI/isTvxl5/tuwvxr1ggqrzGcvCVoiBwJKOMn7KXd9yqZZaQWYH4
3bap7s5/x2R4NSXFYHGKeSw6Xv0iYKKzyfGp3X6zXAmr6xMhwOSKb1m8OI4EsOxRVDB/BjAWHDon
B8+32ZSe6vcOaz4n2nnS95PLhD2JXTYur7kFvUVpxmkMURsjIF8RKQPVH1d9n2gugFpG/R7YwwnF
EJw//FdlaQ/X33y+LSH0StF3Fj74/nwbKBMLNTySPeP9/n3NVmtYLLMmwY9Zj5mDouFqq96GjxTl
tJZXu52mTYxyOPgIByUo6efQ1BFea8ZnIlOptAlRnBToW1jDrY/7HfkYrRca0izMr+tPS2vyKSVM
Hdk8Xpl/0R2r16x2Im4XfZMKOKQ85GZ3AuQXohZLQo1K1Ncr28PVSW0ko8tupo7/PjDi3JszfEuA
BtXe8JT7W5UR9vrJYtqaOfp4y5K+PTxiMoEUR+3oft6xVp2ScpOsM0MjM4Kd3+FW8ACglZHQFrVb
XKKXgv81ZroSuwZHesbxpUapNlLuYUBBFXktalw/y1C+iyV3hz+m98i1v2Wis8ocHBo9e5wjZmd8
o3AKM+Rem8wp93dFLMoKazGmwD2PwHV7hN7drowAGsA7H1w92JJdX4vZJtqiEggQNueYzC0L4mxR
/55tw6gbxvIjvsogExCEFcvHgooiDxyLHLo3C5+YGeXWHEfqsG8Q/6iBQZTJEPDDV6Iq6eJZBYms
Wet10zXIDUR9s7Jv/0KXA7GFEG7HR0QCJjKPARvSyhAjLMwhQRsN8yxZaolN1adjeQSZ/i/cxew6
e7WYFOsNjT+69IX5+MUE+9UZJj3o55gg8b4CcGSGLXRdzap0HE1RSb2p40cAhp7aaeZjMiYmlePL
fGKbaXGedGuq8sa8pdcghotZEZ1hQBicIwf9kJGn6p5LDi0LNGvtmyCnjcUR2mn6cgOsb11Nscq+
uz+t/ZbR8rBHOeH6dnsPPQ8tvMxkRcfBVcNZqXAUHX+uUa7J050bDrY+HZ3PcMnrBvhnFkzulg2u
LE37T1NuhWBFfyrwg3ELw5QCnPBGaDTdB7Cb0X6ElbLx0acUczNt5enD/vcgm3u4vyUZXV3078bN
Lpjc/mWJ5uNIcwzHtboan9ik3ZI1Kum19bsZvZKPe6BZppV+OUbIYNLCgmeasQ0yl6Hn90nPra58
itnQABnFqQnQKbdEcyWUEwwXlDaofG75bRFox93pKSMVmewJJ9UEJE4vGvqsMWpiMLqwjkUD+2q/
dUBrcE0oldUH9oDZvO2l5ZcUjOzDP1UXuCaRT11zvXIWQoyIubKbaruBSv3I8rhvriD69MS5VvMp
oebEomKpNT7JIYEU0hw2kuQV5V5/zQ80Cmsavfng9vkFkCPw8oZNrqlYJjE/0IqESbI/VJVLaGuS
wXCsM8BginPanohkIcSp8kHf0uDzPuWejEq+XZjyT4/FGCeRXQGhL+rwejYqunqLCj98MBWh/ARs
aObWH6WyjjtX3zbsGnVNBxgBJGkaKNNdoN4k1sod8wFYOtJf04C8SUQqU0jSDfySp0BdP+d4I6JC
vcXL1HpGbrtQprQ36/quqAIUv2mQ7lSvfBzkesw7nO2GzQDHIUHIAhUDbrEpfBSU6CsgtpoNgjHC
WhqLrnyd7mO7t9tjXH9jOWQXR+D2Jv9YPK++c2kss29dn90zkrJPp/7GZvIrk4Nx06lrgRP9b/yX
PSc3ZxadWml8UfykM00jMEdxX5fA9dlcFzhEWagsbaHGtBo9aUDyeuL5psvbe0MpthCSwDORxD0r
g3UNIQlteYm3AzLjJTcrcfkTMg8M3vKVivCdSDj5bnbW7kOuYJvy+mvejpBO5lw0A40tFGDufU9l
FNncCD1xw1MjNGChgwZfEEDcBlNud3KEvREK2sJBJ41DHVxG9CjJ7JzWmfsFoRTpPlcLdge9AbI0
RNHnE8va2xVN+3Id89N31o7oDLLzKVSb4SFpuJ0Qq1EYfLwP2AdxMmt3WSyw8ICdFV9redNzzm/H
Hd2k5xUPJEUya5ycDqeNXxQ6k1rIBiUf2pl6wdrFb9Yu3XwJrHHoWPxUD4ihzwUgpUF12MJLBHu0
Gl78ETIZHO6YaKcLh34eLjf5T3WmEWX70F5JMfAKBHOOmTKMrNwU4mbM3cMyNrVwL4PeMyTQVJhG
arMKnMLRT23rvm1bim3RHsjlOgSvZ1+SUWc2J5pfy3ovoiyXcjDRZm5cGL0gz4KFw/vcvu/Tk2nW
+LigBH8O3DiJMvDXA+aRotq8d2u7iNRam6cw8cr59fVaANBTtuYpvMBjNoXw0rCkM+IAa/Bp/EH9
qmubNzOS7l7JK2y06cxKqdeZ1WU8u1mnUGrq1jMbWqMkhl58PWXQg3TflkgJiDEm7Zb+o8Py1okP
7NFHaQRtQXH3F7QpApfgwyDbdDgolsULEGtULVuMxwDDMb8FpNp84Yu2tjH1zPAEfGnvquqWkUfj
vR9Hq3/M8qeaiCdgKy6xdTTY8ckEwMcNuapbCcMBnukep+4vOrhvQd0Oc2aX8ujP5Hr91gxdo7xW
NGJNuNlSuX7qferd1r6FCcMttI5anwPNAI9qoGarinWjN5sJLhf+3OiysJ2VRDetrrBcBV+c+RTA
CTRY3bf9GMZ2DZL3m/eo+aZlgiZkMIBcQyzD5FWdXaxSa9zV9vmiLPoDiqEInlTIWat6j7cRM0UG
TwH8IvGQpLCN7cge9vPp17YeK4FrXKQTtGwXR+YvZ9FdjYLWU3mtIeNVZFV0wLP3CMQmRClJ+qdq
By8a86SZXBkM4aAHuvYhjyld9K8tkSmZ4xwLT5ssOWTXwd+N4kHaDzkZiEsdIM2pPM4Y11WpoNoV
bIBmBjkr8oUF/mUo32eXeY9vxeBVoSfjBB9dSd6lp63oN7U0cLXcLimI65bbTnqi9NpxrJgAnuED
lbCGhQeG0eGf29gHcrURkHvaF1GvmyNX5VvhZOvdFam/dUr75Qc5Gv8gruwVSJgBmjEnY/qngn30
NKDDyRiVspgmqVwgFwuzRvAwQkOt7VA/QAFsYNvwMU4VW1EHaZI1UVNzT7aQIGmCfHo5YR6Mut8o
E2iVjloIk6I93+7aNC/eiejrbEA8xI1Vfcz76K1BGFLxgHTWg5pjafQiI7OXhyERZ5frYLKQm4Wd
seYK6YkHh5U2cHooRLO17BPbNkgllaj2gkULaN8kOZ9bA/hHyG5+ZAcjN7DnBsVNl8EtPZHwNsMU
sZy9BA4t1LCY5DOE3fRmDt66HQSAZJtkOtF0oAUQHGx79qERFE8QYLlwjbaj7h1UxyTaLqhus/E9
U0j8jlcv16JUvO0fpiOHR6gr9c5Pn+sdUqRI+z2XV8DAqjFJJ4yZlsboNj/4T0Fh0QSE5aIi/puU
MqfxI++Tb+QKg9+BGtLBqGUe9H09gPTmSlWeO3NRIn7Ml5eSWd6EIGrUUAGhapK+d4B56HXKGGIf
esir79srgf9sQ40mjfCDhw10gwOI4cyOPtoJ3otNTKpvC5fC241uAdyr2jS1ZA+Yl/ZXKYvRbDb5
N8B+iD5HSRw9ROIsExOUMAEc8c0Q5frWtRxWi40CIsYaBESLC1GVgj3hkCHdRkaXpuXII5FrzCHD
+3mmCV0nYWJ1Q7frvY4jfLK3flCi5RFoNnFPmmvJG4+HKcrK4vmNnPdfRKALy7qYijr8V8Shq1j+
hmT4AZGKYOLmJaaCg8F8fPspZyVO03DaZa/VJEA7gnIZe3vtl7XCk0CnUJ3sho+NKsVOIxYB7o4x
xS50Y2BDiI7sPI5g2TdTGdBUsDf+f3L1qM+d5vzZThOTQOhyU8LKtkJuml7N/83k/vFF063R2ESK
d/Q4lurqH7K8mrLVMsq3DKwXFfFMr7DyycHm6gVnb1+eBlprJ0kZSsWS2Zt0s13z4zluypHGP5XD
Tp6MkUrpvDcMlt2KFgIJfPubZNoTAqduE+hr5cK3xWINXXfRUcHJXMqMBS8ioB5KM99vRHMQpOcT
5lFZ05mHZnsujimo1r+aE8q+u7Z+VHfNU1PA0IU0602HXDhXNaSTPhKNT5R25z3025ZZHOxR2IXn
qGIFfomZY+g4pcLJQb+fGvP6TxqOpVswWs37JAHcHNTADXCxrZjmUexjoo1pq19sK81EeCowKnqo
Xw5QvV2EjbHcaCtNM8R6Avc/P6SEXLrfF4+YKIE5XNtZg7CuF2Rn9DS0DS1AB5Kp6/cIHlGOc52f
2Bj7kJXGoQO8uAQub0b2zu6JHyPPr4hsJXxJTuvvi/06OFcfbeItJ6vxIEfVqYjO8mlKq5qmA9FX
4jyL0T3CLbTAc9c5yvdmUSH3q46n9gqJZN81qWf5YKtaK6J9aOEo2aOlThm9bzw4VEWgv+ALCxlY
WM6sasbJgBpEfafJCDjlhTPSMblpCqr6J7AC0C36XVFMuDAE22FssWbCDd9vRBtzfDFZ8iur/M3B
mzfQh/MS6rAPXbGv686YSAvHox3sW0+ioz6dpXv6plRDiu4K93inzAyUG181bPfGogzPeAiY0MuB
yu2DQgyK881+alfC8YpNhkXNRMufnQ7Y78dZmauBO/CWxfXRLCTYFWXshbrOg7FbTVUqhMYwKgj+
RjYphfKjkeFGu/Y9cF3VXSz84zzhbe/k50AA99h6f140ibBGvMouCuoL4kCE05Dotbn2YmWiQ7/Q
3yGJe8F1wKdEdR+4t4xOFRrlD6uzwYqU4lu09EcRA08Oi9Zngub2gEdYuMlBCC7Y7bAbFWzZLDu9
3G+UWxzNOWOF7F08qMtUN8Z8E1t29sLcPjkhbsqEJRAp1wuaEbMQaOc7UgpiqKgaULSf3sk8UFMG
kx86cU8eQfVaBlP4i7PFHf/TwLfCHdhdz+LbrleaVAs/4Yuz9h/pmBrnYIBM3ou8MKo/h8KGI3pb
GpQmxcnQ5kuzZHjY8NJtlUjBDrWGbZjI6mP5+2AAfYAUtOMPRjacgH0TxUFHSy40hzLHfS0lKBfU
/EmGunz0j6O7fUEF6+Xci0KJrtpNuCkwGo5zBoay3nQfSuzNuYl6Oq/bPM+MRa5KO5GyvIoEB421
EKYRSblZZIQXPHyQnJUWrEbiayXZBr9AksaZxabuNnCLGrtFwWb/x9VSoFGfQYtQUiLzQrfWr8+I
YX5bqaydkIsDT0V/F8He901CiY2ZCe6ZFT4EAi+K54ROCtn1Xdy1hJrX1GtuqPZvrMVpG8wRWdbU
NhadWvsS7VwBM4M4WkMrPFf6Z1w0Gk6mA/L2mCS8c8bghAcXB2Rwg4KMrK2VKK3Ke1lqS7fwg077
k7LAPdVDALw1SFke0zFz6zeiWjOyeVw6doZ29YFFMRhBdFe5ITMwQ+U9PHaKmNSWyguBmD4GgD+i
bBTRN6OiHhLUoWW+kp2Hx8pVSHuK2h6n7eEeIz76ZTt82RiOr8RFg7JVM87mmc+jjszLv6WN+0Wq
5WexV5CwopgxwBSQmelHu5M1d5TC6HAqHvr6bSAOKkXPGUN6q1yhANFeg2nXuiMRzJNlnm08JvlZ
jwKa83LFjVSxU+8WR2UCHfopO3KXPJd/UlmpTonKo+L3wcwJ2gakiiJsEqL6A0B7UGq+QeYpXJSn
lfi2QVFGLjSvOwLEgk7foEFpleq/rWn5u9ToRszbBde2qgQKINx+6mz2kHbTiLdAQcw5Gpdfm5zf
/5zWAOPdP6u4cKt46fJYmKvBYR/zYnWPRo0fpBXrQXEx0TXOLnDh8Yg92AF0oUHIdrRSO5/4Zntw
iE4YTQqH11nQGerjJ2xD4com+7WDb/SdxCsRtBXv6/jWNmlAjv7asZqHkpo/mCgFLe0U8JEembWh
MVtfoqDrc+tNlYb2SDIsS1QYLruD3I6FTjEjhJHRAGBRL2DcA88MqocFXdQTitc1flekGriPR0F5
bKrx4w9fjG7q0yyXGxbpVPZi6xlm66zmO3/JrhUo4c3P08T5B8VzJgmGDfQs5/oPE/1Un8QXVhm7
tso4V7shPxVAvRNd/lgAAdn/4DkVKPzcJNwhkfm77a6ukKl0mgfpHd22gVth97LnqvsV0rtkWNqK
cKfh0sW88OhL5WbFMZXhKubwpwX0KZaJ2GLzktBkG6s3S4guor3FZPBfD6/0lMX0BCM+DUBd85Xj
NSvc03k0Lw+lQpjGeNWH7lWGXXKbtBlt9+vtp0rNOpRojJI9HntNQP1YNFS5RrWSZaEfNxgFUnYi
gkM3XbsIKeI1GH7pL/5uEDcAjmYWUvkO7ZKDSuTQhhhcAzuvaGH7Iw/Qejvyk8DM2hcxIx8uyLEC
mU0Fkk7ocL4qKN0gYjof3nQIVAoKB+q5OcAYn9iW1gLIyQBjSG+RU8qC8fnMXOGDSYxPItdqC3uM
R09JVLhgd5ZxODDEOj7wThugYwC6d7tZA3kWwSdfQRl0T9+9hV8p5z+BzND/txJM7k3FzZlpiWwr
Kk2rurjBZkpT64rt4B9ElbAGbTuvRy+P/ZKGDWjdh6LlCixM7NP1cUa2Ij+8wXkGuBKeo6Wp3Fho
pWsMGvQmT+pH6cMuR+4Ah1GAAZycCfvwF0AGFbFk7NE9S0TOL3aZrNOUGRN+KSJ/z8oijGzzP6lz
35PWtZ0N3WrCiHNDqZ0TIydUT56HKofgWKIIqIO6FGipX7fh11dWW/1/6qZNot4+jnwAdjeSXwJN
7WU5lKtCYp3YBcflWRFiEIprGSsqI34wc+/hoC2iUbntMXxFk7YXkjBRG/Fdaq6KzNsZVuqMAk5A
G5xmZJH23Pg0hVJvX4u9RO+lgRyZITjgT6dqPYdYcNDbarXR9QsZLDVkJaTfEgWp2KB6K/Ae+LBA
bdhwsoLhXAyuW4sT7GJSHT2MhN3lN3uSOMjGU/26US02y6zfCr3NPBKXz4DfN9PZQGST0Vzaz9mu
9/Dg7Oan20E+yDByBaf5QQ3tNlJy6IE4eme+3r9FalyzRYwImiNRQZ7YPo9RjnAp3eQmEeoYAh6r
fpFth0SqG7g99NCalmmcnpBZX8mvCDgelQqzpWf60XXkdYRunVja7PJoS9KmLGPkh1Msye7Ho9Qk
XT0C1dIk4p0rsKkminyNcNKr1P559Y8PsUvX6naFcJGNOMsCmqnRqKz8CB3IC3nMl7EQyxli5zHX
uemE4/Qe3lzqE8Yn3gBpZhp2jfzM+mqMeAbzSDThy36uwY0HatOXtU+6e9m5l6aasi/0VrWmCDc0
IZfzofnDvEHQViQ7+AaqRzHW4uYunaWPJ3CBwoi2bogGxDwV+E5UxNk7NV5JF2C+LZ+8QFHvS2CX
E1pjxBUOOiJ9IhXdNQ8ZLtfXDv+NhURV7thIKE2gK8OBEkG5Zrph+tc1zF/YufuN4hI3n/YtM3Dq
3lX4Y94OloY6elcRI7sFhpYViJ1huQs7DNm8QoQ0xerzVNmtx+J4TaiqEv2jBFu4o/2v8POdID17
E0qCPqHIr4qgyg19QSRqbfTs00anhBb/gaRJIq26vfu6gKDNSjXYq1F4Scji5+62eBNBIKjYUMBd
E35JLVg2TJ42AeMS0a2PMCsraMEe5hdZkUAwmaS21rIuj4m2giK1DMPAcQBbmM9ypvri++f/3pdn
t7EBsliF7mTZ1zLRvuP5OrCJX6rS/DBZpVdsNQO2p+VyxVsmH4aAHEzMGA2Fb2YqoLr/r86qIE0d
rsXfH8iP8Wg/g1duaqEP1t/QfHS2z8n9ooHTrW+R9116RUD6XOq7eUf9lJAqoROAB87OqyLVak4z
uvW/DCiL9qXKfe1FOGiWj7/PWMvmJtA9umJI1SYsLu0fVyK5lmqg928gaTJiKTNj8zpOLvgxanqg
5qQQBHgc3khcVeZ7Onco/tdMIwIwfKFj1pD0DJhNauCDczr49PsTdnBXhUT+Csjla9oKhT8F0nia
OIChPxQNx/VlrQXkZWFylkBwK6DW+7nqQkleKAG9pyJpsC6lzv+YJXxij5gqqyRpyG0I2fxvL0Fq
foOVmjlxUzLAXS1JUJkI9sNdRFstVHR4OcaXwY2rtUMy02F0TmGpvCqTUGD3uGweAq2oPE0bs3JN
wwmrrNSmYlucxdEkp7SYtl6D1IPJZrE/IrkQP7F4GbWhuUDfKT7mLxEQaxhJP3S/MkZPsdKAM5CC
gT6Huf8gEsMv0tJo6Ll28gC87cVLhpofkoHbkzx2hDvmDoxbOoj5VFkmg+a+b0cVQ6FOrXKHNoZY
tUuQwALZAgHpsNaA1pQFfkAIvQiwJyxJchXpANu03akQfA0IIvaba1lwpqpz7EqF9j6n7r+sTYYs
BMtPAGgJunnF5U6xPWB2BJo0R3ZHpd7cARFJQcjWDBqWPb9lcSTtFiz6fekTvkRvjDtO4i9gGJpq
+GobDIlPZB79CdS19jNXfu3spE2GWv8U0GVqG4CDbgklvPXm3xRZfeeNoKrtgScqirl1+ztW7S6t
5rdIJVuGSKoj/xJBP0iszIsWKBzSAoHQIPfd8QtJjEGuEp77PUA3w+b7AGyl8a6efPkaMv83TieG
cEJGFID/h21+iVWegvhf9boFVV+pOtPiBEyJo4pNq37pTYpgb34lWDgXCALSJOf51gB3VycKRpUp
g/NrbjDN0fw6FCLvJvwFR88icmGqKwKmNS9y2ef6qNQf22kIvEqh9jxis75C5a/7T8PVeV4JW4ux
Z/C3Fxc/ybPmswU9bHdHJUrcXSheTPMVgmVgQZ8Q/Wpj9kLDXB/c0OLPShuPZQTVokbbfyXyOLgh
mw3pe3kw6GsHDALTBP6crrsVUDKOlxXjBNpA/8ru6mvGuCvvf4/sth/tF7G4O/iXDhmZvf3riyj2
TbAVecpiDmDuvNbkFuCuzkdSerG4g2oY7+yl9r4ulrAaQn5TkQfXLgIJNXnvzmS+MNW1bmNLIR8y
umsFUhqKS6j+sIAvM3IF678ZOMQjJ+i0xHbhdLFarqreEI3drz6jxMH2W5EZpp0P3DrIr7kpnfei
pmDIaui13Ag4h+iQSNQQUC4gjwpwblQoZoheaIBnD99KjKIa8wi4vDyemjlfWbJRvWRNgHL2eWF8
X26qGVQAmd+vTfGF0EyQbOx1o72bkgPtft0n6cQPAWNVOTGBrqOfSyhQadYI5ilJLivomhn43nGG
p37AthKFWeTzm+NtvQUPocrfVlZIevmir7Mg7RsG8gmNyGsKtXgS2HC9ZCRSvHpuJWd9frImngEK
ssEfacSnhwj4teEtw8ntheT6xVkL0r9USz6tSq7ZPLAqQsaE+G+gLG/C27w0HkxNdJCYQ0azQTt/
0+M/gzkgyAEp8/0bsSOLFeSYZUFmx0uEM8vBJ8GS2uuKadayVVw4EZR8tUv/TaZ6nDR4cFU5dAb4
2amMPeIIot+vUR+ICeuMYe5+Fp2odQELv1tbB9M7ufU6oJOaX0g7VNLEgU1zpHG63ycBhtBhb1x8
mm94z7qN2qZ5T13t/Y65ecqGyIOV3Zq1GxqQjpGE4cFtyoSNLocqTPTIHE/KuJP2RyT3ZgFZdaiF
BkXVQZcjyKGGIMtMaMvUntbTFVm5rWakcNsIetpKdMvMuAjRi48LCRBYGyb+D+ZNml+eAMydcuAD
CvcSXddQWauzOlTlxA35YYywlnOqkk/iDRtxNfGLbgvHvJ4ubolPrCx6TEWZSBW4NjhTNgEY1tPl
8HRJ9vv0f9Z8VDBsEKi+QFZVgFzakjnF+SdmcVUcjq/dRekfxc3yUpMZH4Bn4518Qb4anWNvNGDK
SKhZdrraXMV0rfDAYKVP07W77tkS1ynD0c5556nsV6Xq/g14q3BO18I95lMMitY8yic6mEtKZ3r1
cHLBq0G9Ldg0lXeXL62QVhaHlBNSayES45B8//HaCTWh3ofZPCXeMp47PFXnCGOXlHvxiHMky80r
zwEKGMuIgLx4hk7l9ZGd4GwAMy+ApqcTi5vj1csVa+o3wknf1MFO1BjVpT4DxvdZzZ2fEr49u2J7
MRmK/uEVE1npw2lFQK97vMQ1Vo7uD4u28o25A1Hj62Ze6P9eal/IY9v/QJjRIWOpLGFNUqK442LS
Zfxs2YMd7W3OI0KwugKowUqHqkxKvlvQ57y24UEh0MG7a1bGhZd8K6duv9/JCR02Sb9WtinxOXnm
BywCC6U1YstY5zQNIF3t55BxgJhSzjLV/dGBwlIHQwUATI+Y9pQDy+hdkR3UkWKD72kvcP4WQEAt
K0ONvGvgbyRppCVyK5le2o7aMwPv205wg/XyyUdjmse0FTlVUQJOeDWPHq/WuO5ndKMOFUhhQP6E
amDAubovmRxuuDy/SIdZi+VjuwzlIAGI1B8XC0uJ++xevGE9LaIx4W3UPqPznArswWxM09cx5Iqe
Xt6eE/mZuCQ1iJrf9exH7WTyxMml12B4VCj1elrn98C2kezMGMqIDCQDGiwFKZkpRHjFp3oRGl+9
c3cHkg27UcWdUiExV6iocbERkK06ReQDA2C5y3VQTPNjou1igw/MqkvQvq8ucn9faB+QIKOD2tYr
oyDZ2L+elBX4iMLp6VQUhjEL5uw0tl9/VzkInFdv0zO8wh4CRfyarUA8fNtR80yEVG/FP1CebE1Y
u6Cvx57FFOBrv64G3AWXExqd+1+rGOmqRnrqgbTNfzAxGkivicsI5/7iLkHaA0J7jS/r4wnFdpk3
UPsK5KaTzCJYuIEf+pYYXR7oPtbaj+Mp1irGABzPwx5rBLr3zApaeuPQAfheUNNXKOu0RSUc6bKr
VE8mD0MG1+PfXRaT1YDdHRA2tiBczJvFPfQxPiKk37/kxRezhNw0MMW3VHo8oYdyocXqwsd5m6OY
Yo2EXx3CsgGY8tWvOd+Bk3JJjgkqLi4D7F2Z9jwxaLAwZTWc5pjGlwnIUBEwjIxu00MJvbLzZuAy
zrUHLFtczkIymer2/zw+WXzowDAazyW1srGq8Zh6rNNyf1JgtOG21vMAnM+ZTVoNVj3u8c1KMzez
S4jmyjiMfq+NVwh/MPOL0yMd4K3O/A2zzFEhOWCYNsIB+42TBOYQ0AL1wIsSwt3Pe8I7wvHbcwLB
DtuFuqiXn9y8XjiC0g0MzE6OXF0dZsjMDmLKcKuFRvMPAiGBvp7ZxPgoh2bWKe9cZcdg8avJ4Gop
Z66XaGcPoGkiNqdMKbr6mUOZQKlStGEbMTxJyE8GKD1vPk87h9bAFJV1gFHgIieK3+Ye7PK8w3Q/
GakBo4RwkPQ8Q9PVq/ECotbQsJ9fMgRGyUQjmxQ12LYb61Y60D7valouas9In9+YH+VPtidvxc1i
gF6CbHSvYl7yb7RdZcBqosDUUO8yGFHVXZCKpz9OiVJUFSks25xPwxuk3CHhEhDq2jFTf11PST3d
Ft35p7gqqMAuZN6wNn/HHQnLnnd24hLnZdALwPQBF/aITRugpHPAp9pBpPz8H2c9hpqUBmOttNA7
FEGisSl1Jkc0wuIQJsF5wK7rwFZpRVEGppTvAM2qB2tknF7UIvD0UJhnRncT1toH2c3xBwOQQyOb
tijlUw7uywbj9TKaFVlgpGGXvzR753BI8uATyi7gT3HAhMmFGZYY63eM7lZK4Q8sXbVEx7V/SiGD
7DC+QC/wmNrJSBwtmg0Ndc6/UEGzgEpy1KdCfArFkoB+fTT1aNk7iePrRcSTMOKxZ93nwliLOEx7
nSK+vrae1EQwpEsH5tuDQzoBVm5eZj5ihuedIsHnZIObqiaV72dxihXlYbYuPH1D683hj+NdkTT+
bCt9osQQVRy6g0Itorvd1EC/wyJlhQ4P4ne0oA4NeEEIyqmOk2phG18JiDkRUDQZYm5naN1ReFXs
lS9YoV9D55XyA3PuZmTQBE+Dj6OMApqB+NID93Hae6fmPRfKGQQd76qd7mC49Vy/+vxOFpneZ9LL
kl/CYFcVTQaCEZdjaKsI8UxQVJAzqST7Jl+lu5vP7VQLUaL5jm1rQzuYk0oebngB52F02gRdlHOh
WH3bw1AGiHGnJx0xVPmW4q5yDUsCAoG0Jv0ySxhl/3nQ7FdKSzJLVbwb0gcFYSBABy/z/DJZuUaP
3WirHKYTxZR7+/8/D49Bw7BwKagFB7DaFjfzwAnXlKXuwcXooHuH4jeRqkuQXEcSTT9xQtNCE10o
XTaiu+qH7CqS6+L4bkUV+M4N4MLa0vCcAjEHIrCoeKgsYImOMRyc/VHQlEM9M5c27jZ2Mp4dnObF
zEKpkHS9nFrfAY5samISKbYxb2hDIK1u2tO7yKaEmtQ35AwWHFjG66JxIfa220kp5BC7cD3OSC2b
8avcyaN4qDeF3s5m/z/yMqD+Eebtop3D+RpUrIeYTb+IHF7v6kIx0d56PQ8IUNZbKCytncERDyBc
YxNXD8SeEWBSqE839k59I2Rb6sL5T4NRSHqRW0U9pWEOOMVnFc2/R3mqp7rec9oKYr/Y1zvNKT4/
qoTLvl8DGcef2LrWo3rgmU2J1O3q/SLu9n5stUoPJ2ELPj3eRa7KDIFQMU9hObXdYOJfPkGpR1J/
fsswkqHOrPN/j4Kjr9Ndns6v8D+B7Ag3dGapJJlocfmtyG08nc+OEDK8LccaAdB4bFqVe80lKsY+
rYY0mLG5tzjZIen1c+gt2ox5cvlk/a4Z2ZjyawsVaRyS4K+sb2wih8x/Je5IfU5hCb4vD4bIjJ3b
U2hSJQX2/WkBCFqskcj4lNY7/IwsAsE92oJIy91xK/yQVaAXX7TvBB27PtdSnIk42a1LnV5dBEMt
WcXzYF638ISCLnVkmqc0MZyoHL/yAiekQxxJyNsqQiKzr+jLOFJNS7QIcJZdI9Mxln6QzrriT0ZW
GPwoK7oNtB+gXixWpaaY87EiVOS/t3Z4nEg5kMdjRP5jg7JZtLkR9LOvpo6iewFKYC5EX2oFh4n8
Q79cLc9LdJ2a1mgMc7HC2voQXpBhvRmb9gKi+PORPtj/vlU/cYpQ3vT/QhqaxYiu7S20mRsN10gr
syw28k9+y5yd/y1OCehd+s9nJ+L9QGk2dIT6uBiXIRAAAnMzi998e3nSSDzWUecRnd8JnH8326eO
OOxZMlF0uELet6trupN6ETyuAEq2kWGmI5VnIWs866EZ3E3PJW6KF8xL9/WsMbSpvWcIFNRlPYLm
t4HyhocQQr4VOw6ToeULB1QmzP6xIluKKfnOhzVzcdBNH1xbrSE+ijRJ4KSoWkI3SzDWax+hPfsy
UkXzUNrqGybBFcnTuJm+DC94Pss08AbbSCU9+rE/S/XfhaprFyFwYxBLDKoLeqjJV3ukD6OLHuUL
K/L1PyxfgI2TUR8LIF7VzYMupwQaY1bZLW8T+AsGUbmI+xV8KFIE7jeG1kIs1xyApbuDWrE96eWF
1jvVhy4/6j8TVlKDkkCCd7ZcSM+5pXgx2G8B6G4nxRncYxTDoFjTEfwye5GWD4SbcffZg8wv6nL5
lC843G/JoXXJJ0SZ6+I0OL9hQm10FPeLnBHHI4whHswAYgchoS0i4dEawLGHMPNTK9GAxUJgl/IZ
+A6fxve165g5bBUVYSXBbMAhGsGI0VT/IrmHK866tvyoJ7QkeKxMjQa7jle2JGpydSlEW+Y/DZ8O
5rdqeFZF17Cl+YhBH0wFxqEw2f58unSIRVxBzN1WZ8Rj3TOssYx0u6FMj22JZHilvkHKeYPiXIIP
ccYBc+EL6iLUXlAuD1L7tGkzRU44cPu01p4N1p0cE1cmpEgo2D2NVMfWFiOganDw3T5naM4wIsXD
gCTcILvWaLHZPC51j3GHBZtJ54sQMQbeFypFmeu3BaSuLfjQJccujo7wnGuUvY4YxaCGtSvCT+D8
EfE9HPUDDm8f8E5UL0LPYbMZLZWsChgKtxUzgmi2OKYfVyDyg2Nyh5uUCSuszXoMYjq5JKRcgwjc
KsFx5GQEbY8p5AcAGzyKIRyx2RcffMroEI2fpDbLLJXoTU+E8nWPH2vohOfazOe9PXkKNKy3T1hy
iwuJ+0OS0TgtDtqDs1BZWXR+CeMd/Ij1LpX60G502ySNJxKhP3Z5mYywjgEt/pbV6T8HFOVhNHUD
Cn9XwnxnVxsnuaZbgiR/v94Vb8ge12MDm2vB3wL2HGUUMDmg9D6lCy2bKxpTYD/l6E/Zwgqs1eVM
4EmDIjxDARo3VqZsaY9m/VmukH/elJ97mo4zvyi7zH+7w9jkTV1bBx43qCI5RPyFc+L1FYjDGbnu
GcyFkTAdgXwLqnHkPDsoeKG2L7qTdM/RW+4c1mN2QlFpLp3OG5JWQffqYfSUh8peC29LQfFC/Pul
BFKOoEUsTn5Ds+Zf+vWpppNygOSVMCP5s+d9zMkbUJ2BphAeJURCHoi7Ln2Wq2vLYJW+8QVqeTR/
Wlk36l1VrCgoyQi3nWeOEA9QsbtwON6R4sJAFp6Wfspa22nRRFQPeLDCg1bnSxcOPzgPa9FkgnRs
z1YbFlz4pa2Sec/Xh+UUHVDKA9nU1EyqnzyBerwz67IowIukJUCqVt2ZB3kgTwHOER9sJi7pwsDx
uxZnd2c+W12ubx28IoHLnOgmG+1WrMF2gvrv/shIs0KZkaRJaBEPF/jT8hHaWyvV4vhLyytJCeuP
OCISQTY+1y+jsqJr4cBv32K4dgZ0yVyFllD49l0EhMipyJkCchMiEtKGBZkdnhr+VMg5chtIVNK+
IBZYpwwUxqUP6SronRjuvobn/hNougTRZH+0jnw1q7/YT/hRXt4Omr9vU4MUFd3aN3P0wh2p59Lu
0UeZ7kUosPMGfsDGtR4y7q8u5gEvM94KklsJzp9r7ToEJtU0f6MHguT4AG2n13lhmTzGsvxkm4p3
ODeSZ3tdMZn+bkfZlcMxf2uCkPfzEmgRGLtInp0E5/YkByiNB/nBCHscrXIgGxHgSOvl2DfW+grg
VM4E009KicQCmRVyOooSk8WkS+Fd4ANTTec2tHd0tOlqMKTQnx+szJx+s3WXi8ZU/HFe5SSIjh62
X1fo9x/GXjH6ZcUh+pWkUmxY1l/2YlvI5o0YrLIufUaEqXrOX9P5/PwFpMvvNVRYI45oVVbHlNVm
twmTGrKBkJHXUgarPeTXsvMBGKDFfAHA+5iwnRd/yLXJ6pJM6PVe9SwjREh61sVVBEjH77/pllw/
Kp1RNtDQB5t23OhbPcTkJpugBV6I0uhyuifaF1oDZwqsU3F+KQGw5H+IWz+C+SG35iJNUa1n9Vx9
3IlTomiEpXs5ToEpbR2C9fxdYKVkPpj0DXV3ztCO7UF55z4naJQEyOn3J1dWF/aDC2BO6Tva0xyS
qNQuJHeVkOl/3g3Ev2gsLx7HMihCHzA5A5voP7H5dKQHPcSZ/EPrgY1+mxnWyh8N0wss3druiJwB
f5qOjJUot7CxnaopxD9+INfQfOSSyjT5ReNWGNSlgbhf8O7kxNFsTPdsI9fPmRYlbXltt+XQJgen
xE8SC0FW4LzHgWmoiCXZLHAXaWwe+1j7nJCPeAFwKTFFdU40Uyht+Ox9JwXmeVM2LntrlvYkdJcN
tf/lWKyrQH38veAB8B4tauT/VhfGRgdfhIdA1EGBNOezei7A12dClsjLSmInyXNDK+B4UmnUjIyk
3YdoIcBTGCzzG51XGmBi8ps7z1vj9yqEmd5TeQrS6iZgUlTHYFvilrTl8UyvjZZ21fCBZ43kiA2J
aNKUNd1KdBrghIveCLFWXGnXsI1nI/upiooxfKzsD5FAxECKVJ8Crq1UZ59yvtEwONZIjSKELGe6
fuCjJw824qK5wugV7H+07GeW19l2TBxMOL0mcjcoAhq5xoKnYt0qAG3sxmSFuAPV3bZB57a3MAP6
yMrdZGeYiDOPvJ/cySq67ZxTfyqtiBnXncG3KdO19dUGTS2BNsN24Xrm8ACsEl07q6sSQTuAB7UO
nNYuJcFXNmycDztlrvnuHP7yYM8CKOEdI7kosFP2MYJLDXJadlh+h8Mm1AYsLXfxztC3l/RFb1Dh
Kk7yqsTQQ7xAo3/URonkpOr72x5L3SoZO4wKBNCZA1V0Acv+lkckNlo+N/pj6HbEzjO5/K8TX5cA
K6tyPsWIwiEmviEjb+4VlWeH9Jr33tJTHUnVk1wssgxzGCli515xqxH0D68kf8JOm7T2vOKUTHBc
m+YnIlo5ds+IWgB2HieECnGZ+HtSnMZ6wHo5fumqmJqUwovcnl6MWcebqfa1Xab4W2fcaK9CzWam
9wAxgeW7CDu43OfK3nw9+e7gO9c2nWtIQ93PiVKgsaHiINjenEY8aK4CSqq880EYbEAzr73ZBjAD
FoDV0A6HlIwnNtHZkblhcsQK5uejv13y7N1fZeYH6LDFvC4F0g2EUld0pRdIzC1G6gUvPDIUjxIJ
chs8J4DTY2+aBKLCwpZk50+AxYceZLFsQOJ73Ph0Y6skJMzj2KTM8hXEBvmbmGkNAAKjWKHcaq6N
5lsKmn02znE1iz3VLt856ZLiFZ1eyR71S3M8lQg1QVH6WfDlGH9sxB1k7LSobbG2ZIwCi387cUlC
Th8Dxav6Iya3cf/CIjQmKonenrM7H526Bps/Sz6l39qYYbmNeHI6WhbggRktEKyx6dkvEGYsW27g
bfSpPagHN4i3C9/XidBEDS7zeWrLHhYHaP3meViX42ADVO6R52aJ3zkK4aDzn9UjD+Lh3SjRLkvM
msuYNDFA/f8mcjyM0ZAupfM+/3ziSackx82VDoSiLoSCkftObRS1lBHJeHCxhNv74ygTH/dNYzgr
yG/cS+cVAFDkie0Nq9FCnVNIPn2omaDagwsc6RF+WU65/VHTCcLDNgn+AkOohhSfMnKkqJ3goZRC
w0bWnbrP54UAfAlnN7X35euopKhhCtXPqHaO6pXG/in9xomPSiGXyJ9qeA28TfqXWbFESYacE/Cm
aEDb2zKdtduTv+OuZ5SmwpjSc4Ygy8pd+ybkqlmW4SBhXaWw81DOzQwEAauLzjYUpFhtgtXNekFQ
QCZhuxcV0Y03mnvyM4+v/Hx0hgW3QuGAiSP+BZJKjwR74wgGjPcvnOpEe/QwOixa0YmWphw9Pij2
qw3e91udnVMfeWCXRkXSgtW/Qkkt6gYEDWfh3+w2knBceqIdAHJ95877WT2qyHDBCzFlyDtUkz6d
01FjgbCeJ/RsFusSvD0/xQTf649MRLMuIllYTbLUkO259T3rteNHdGYQFmVEQy2eXSEleewrBdLM
ATdWjwuR1jGCNrdArotl1jbeuhgW+O5sC9dBNlpkh/m65Cf4ye7o7yPUhylpbkX5ikjfy3OzGZGB
IyONX25j8Btt5T8pDYsh1+6uAhoMsjLpTZqx9+bYMLz/0qZu2g8ikd6ZMzzqu17hFiNAxGBdwseB
6ER+AnYIVJ2gJ8AFrp1RrWYmq7XHCgOo6NTqeqcKHbvdeLfJHRIfJcYaH/E+gaTKyEUQ/4YT75bY
Mk2U0LNo+yA1Mqf0X24X11cVppaKXN4gUKBZrJ+y0xN4QIQNoXZ3sgfh+V6+Isx3tT9sdit7AIzR
rrlKoOcssHTeq8XmHInyEqwVDEhn2DZm0f1fJ+gQpHQxA+Kd0J3Jn+YHGDZCNvcbTFICoeTp+Jxy
KCtSwByNL5hCL4qYh39gZNF4qjFTcKRbZIrFkJuDdSHYAajjC7XCe8esQR6m5nfuoLrgtfHlBx9v
Nf1VkpQGTayGVkri7DMlzlZoCMsg+ES/pIWuieupOjWlXo9wfSyd4gm1ZasOo7KPJzbUqeJ6fQIR
ctCjnm7kfXUwR3wifwjDnTyJx36oDi2fmRbk2GCSFmI1h391FY4f5ofSUttdGlpnZ7/rQaLZDHJR
pIA+ueSTvzN6DeeQ6P1vU1VWbz5/QO5q7rUozErZOFeZLpzQ1H80VndKNdSJ7SI4m6dDdWGRGzBq
BpUIb28FKvECEwWkei+OInbzakAEug9WMg8qfCyQV0JEP3nAVdUtlTFEWIWr4unpWx6XOZnSWb7k
9hEE66xiMcVd8xCpMaCA1mpJbqlYW9pYWsCbjCJHAQzFBHexFxDTOL7BUVuotjwCYmoIOt/jggMW
1CJ1egPNmQBvRlf63i3VK2WecOOBBfmz1ms4KLPHGCv23+U6/cOq8bymTk7F1Qyv3TNIKGzeg8rX
NakP6gm2etR/8Yr7o5Zy3sRhWLT3phrGpyosAsSkpszrDNuiCLEowe9N2g6kAa/F55tbrHa72g9y
vLXslW15bgUFT40ku/oHXxzIvKIPql9kLid/+WWZE7OmNeFGLvoPZEpvL11USgp35GZ8D5r3a/I9
W/QUJdkdN9NWcOBS1pFuU6hJUemJv2URRcXv9y6F+HszgeF1eKNlZF6d1/lGX9HUYP9WqFAtrpwI
jjCb2oGxSGi/Rg7vknXKP1C9PCK8zpuLwYe1OFUZgeE8HEHR2GP7ge+B2RAEqHXl85yf+Cxe3ZQH
BPo7cTVjeY9KQ4fyA+JSZ9XvjT10RL33X6ZDUSRYFNaW2L7wkU5NhV/PoJvxf1EP2dYtFL63aYOQ
1xqCvFE9RJzviHDgqevaxOZ++3m6BYMLQODloPV7gfI5BHjqkEqeBOdIlPPu4RCniY+SfdfTq8Sk
TCyNfLRhHjFQRGPa6Tq3nGPFZ1+W4v9IQ64VMxC7rOEL+w1HC82CzFitztT/JCquHOss6tdcuZjY
kdfrVd6W57S2bSdm9SEQGXCgl2joTHODI/BjXP8cB4eNtagKZfgRQ7Zc68qfEhm/NFC8QK9iqTMK
BR/Ys0zpZC0k07cc+7AanhX1QvqnIwChZFpN0ts7GQox5+KxGkghu7zBmuaTZyiLQm6myewrcTVV
Qo5lnU2m+vt2hH1oUwc5irOLnI8p/NdGs+ASz5n4Uum4qRGXfqE7b4JiHfSvew+kinI/9qDciNhq
pfnarsJFujyQSMH6XH8b1yMMDpLqDPXH3r/Ozh5tYdudNr7wx9FK2EU1vOmYHv+nbFvBeYP2v6Oa
cq1a1k6J9n9VHEg21u8zfWNiMgX/v+54ZMf8QB8O9tmmZW1KSwAHrn/4Ri6QxFjK0p7m9638Cgyt
56vtwgr/Vy0dER/rVGMO4xX5T4ISH9qOqR8pRxfGqXUDRC/xaEJ5Uucn5EpxsoqQlQlNxNGktfDD
ITnnF/YNqMp61GiOvuMCLmWfi29XMQZpfyY6uCxk7xdN5zvWiYk/rOJbgfxQO4TNerVDVsZhYRQm
tNDabDscCS1RQs2b2/3BN1a7K7QQQ03J1Zxdnpx5E0FghKHrGtOp5R9aZbNueRPzsKaPtc8+RSXS
tkrMzw9iTZRzdCk3WhSCt9HdLMp487oSHFXdN/V4Dv66Sn37jn/xRcaNNyPGJwOZ04KsQigUEc8L
B8kymeWYnDG36ap5L+WT3l9QVmOic2zz2VWPRt4X4uuk6ktU0WnNqAa7nFs3gV7uk/zIbiPlg+yr
2v9EMDOf7Nbo9jYJODjJbgIyWUPMjBDljlBc3quUaoOXewzAxq1fHghgZKs5/6U4pMhTETZmPI2v
xnZ+1rMMkuK+TvlTtRqlcBjJuHlCCK5/ceg052p7+kr5FH+bigUoyScxVh90FU/Ge3CbGmvo6nO/
D4iK+y11oQDul1q/xMLjYFTqyOHlXxXTdZAwS5jZWCO5tTiN4SXH0/km9gI2gX51CT7ootNpJw7x
hOkgQH4PyjQgD9EmgI+5bH99faZ95TmuRRJwXmpA9HMCZ3yLvPuA/gmUWaDBO82RKfL45V6hr6nk
BDHouGwVjr3tfzWTtxhEVRbzuRIAEIAY/2gG1ieUDQn0Qm4GsBMEItnXyUE4m6yf1BfPdMb25KJL
RcF0O3wBjHziIrz0vsmRhjWG5F7VxpA3HbTm08XngXXcYUWVkpeuDLGX8i4LMiq1dNXfL5WVrnE5
rPXx7qBqzRqXB8xrNRxubzFEgNqfu1j0sATEa8tDTt9+ShAQh+hUnodaIZJ+rU9+t40jJS5NrO2b
Hh2yWk/K89D3Ge0qli8JNjNv30h+z/e/GsTH6j0BEfu7F6vlSPJqNRBg3UUeLFEIX95WdvYReZ0l
LUWd337cegu1e0cUu1kWm0EA9RZO4f49mUCb2an7j5YwXqkMQ7Ckrf9qOdvvY/Aufgtfdf5byh+b
L3HSCwDTE2q3R4hy/aCl59pqJa4JEKO5xwiuMUKRQ1tEH6ZgVzTQUkN43IA96jeo+JictArzZJT/
lafBwGBoZu822+XoL26C2cPSVqFuHaGQFiY2AzIzuJmfWQ3uwz4A4CIasyFhBAw3KdomhBJRh5Wz
xJN2K4UDr/oAme1AjEDqdfygqu7Ji5Uph3+gHKxJOZ80z6M4zPgtwimtDZgKbb+oNLAb5BVhyG//
4LJNFbwQDtJa5djXxA1NM3vpRHDJns/q4KeoHBHtygPT0Nr+lAbJMhgIczeTVkkPcPQHZR2M79v+
BEXJdMJKmsKUs6NRnom/OzUtOLcl11V5GXNNmELXqmtMrYLaWK6RaXx/LB5bokzM0zVScbfJNnzX
PpnkVNOo3Q8I6YDyP6giwg+9umcvS9FIYeDBZSiJ788KDvTGc2CpdNF7rWzf8t9ujgGzsTmdrnnV
e6X4OdXspz4zT2eESvGBwEhMjsF/uJrASdhEhCPXw26cWPVNhXkTglkjMmwTCQXWae62PgKb7ZvQ
wVd3fRm9SNx3AFfBYBZyC8eT/euBDx8iNPLNgSvxmtpu1+n50T4sCXf6QD+OreAxZeCMrRSwmkoQ
PJem52RmL+xQeLaTsVgyWB2NCgLrC/7xtugjc7DmIADJv4vCaibVBhif5LpXstqt3VcGXEgkjQLy
ljjGa4iuh35Q0FeZO6OcOktim92wfdZCb3SSbSw2xwI55oV2TfsE9Qn/MlDx1B/2OsXHHcYqB2G6
Btxkj++xDZodA4MIg6qbs4822G1gdd+DJHN02KjnBQS3jX3EAjLQEWngJkiX6iqru/LKznjOXNZL
y8jKU3Crz0lLnWJ8h7on9hYZhw3+34TzzrK5kJz+n+pyfUToxzkjov4+k+Y2tCl2laNdB9pTHzCl
BM7p+71W4FSM1dDoj8gXFcVvmqZ44un9GBqF+7QTFd0VvSigfZdfGvyDJYzByZC9fpL529dZmyKP
6iuBjkpxgSJHH0GTE81oUMzxb87srVYoWu/XdTGzbJ+I44yuSV4cZ4UcdKF96Z8IS8/Gt1GIigWg
qIAOhJE3SIiyYWDfmUOYm+ufMN7MVfcmAeCCrJPH0QllGzUHWS8a2laUd3oQrFS3dXL4grSu3o1s
Rvr/XGvy1pKaz52p8qS1OpZ0UQ9ibTT7lR9O2BMHU1XRw7Q8uXSrfq0f/eZo8b63TLGSa51XlnO7
GW5p+Q9r+mz/80imGv/WNATgVJOjOryit0r9fMxwX8saQa9+9Qt99FPlUQISi+UwWrPbAgZvgRac
TmyDs3bNILuLSBpBQchQRtv1BR2moye1MzpUrZe/WVQxmwqZVSdvfQMZBJr4k62vu/aaqEbqYXaW
smwOJRwg7YSqBrF+wqE/L8q0FlIwfb2OOACLdP2tV1PtFpuqmlpeGvY1ucW/mBoPPnJ7IfNjkSFw
8Dbuu1c6hLjcoKjV+x1ZAvbFUcp/SqgfGuYSD8IFxFPR1QJ07yXGJ6Ek0tqIQBiH5+fBlXGCNWoK
gBPEIiu1iLkLwotfWbPSdGoIdBX3uEWhS0bQRzbsaGhNTdhEOLtRy41UbjL9IbeeMtl4FvDHeoMB
sMWvr19+dGiM8U6EABzFz2COn0vyDpGw/xu/t3t5MMSmf6Jzzs+ptQN55RP/ewjm4wUnoAXYDtZi
LFivZHYEB/llgkYOttbTAAr5bfeiHa59gXspK99UJT8Tf6YrRO5x8BPD7PPaCk58vEnjPIjIK0kM
VjVNFf1sT6jR/+DdM/TEbcIEF4pKCXr0VlXpw12KkUrNkAbusDwacY9SzfOnSue6itjPZB/zie71
wlYepZpuS0k5A8ptW1ouDAD8SNghwuI/9jrV9B4G+5h9JkHhyvqq7q/escWmdF9k3IbeHSWgUCFp
eIarl01SgvpUT8WzWEqDWtf+f502UnnnE+OIxFiZL1JxaOZKWqvGszLRA6Xiqk2tbLxysiW9uH4/
9bzgkoG4I71qbLW7NsB7RkmER83cggaDdFbk24k44GDT+l6wAYUxe3YnOCJAg+9MX7XalCpVBLg4
wS+r9wNrzirN1gANi98F5oxaZsOINeLCB8CCcuZ2Wgzr5erjDPYBiePuF64pdzrK3y0D2swgYtri
1Lr1L8nU3rYgKBh14lcVTh2QPGOqvHDw3TyxVbIHPKG+ajEW73u6XSS8jQW5wE2bTYKeAnqG+now
67QjX/OJSFe4g2S3UjePC1ts7/SU6/OlyUOrX/GmX8qT5n5EqWERd3/nE6VdeNMWLy54rKzEcVIC
D9ReimMjkO71H7yg6wpHbwHnMaVgFlGXHaUMzAYr0BidsajAjBmMUIMbh4Eld89f9BCIAXYmnQ4I
Lxjlxq/1POQM5jB7cc0YjJvdNTP8ccVIWMZSI5XO3ey36bBCMXVBLBMmBGEJQrZ78mvJXO08OlFq
XSB9e7ygvniCLLpdu3VhCi8cj/ucenvEvZkRyoHTV2Bdy01RY80IqmL6qYIIVEZxBi3N93UUFHn+
iVALxQB2ShnotOFOqgBUcrlpro87x0XFTucNaCBPIQwL9hK/wuMzAQ+TK0bj0q5NCp+Lfv+e+VB+
aOCqBKMmF6BC6pfhsteWy1/adccpB2aLVw5FS+JC+jATeWWXI8QyBRLkuzXzwkaQ+NeuSlfVf0UR
HMv8sHSQBM28PCLJ6XGn+4ahXAGYmoww78QhqNJikA8tZSBBEVOEu2FZR4WqgRjLlTLsfGUbH7Te
MzlaydQwRhIHqqNOv9A1Jvn5GmP/tQDaNtB2ggSWabYP/6DAaJkR4VRfk58F9YADGuhqjXk/9wZz
KWKhOWgaKvlh4loIvH0zjAQ5tu3nIHxLGNgEEqalP7U2k/G6SBKTl0uZxf0xblShj70rA+bEurbP
tuIoUMx9/+/na7Nc5MbRcuoOp55SiEZ/zIiRX6QlPydaAPqcvt8B9IGClLJlXce+b9+cDucEIrjs
bgn5xsamw6QYqRCi7mY2rir5veWai7PC+T77uoBwjLJQnbhYxkfy5KkUfhlQjBAS77yq5TcS4xkl
FThYpKEkZ4w16NDycV++5A8QEsXP2y7XKdcfXrecVLjtB6sOdtkK+TJ0HJJwjPfnHIfICCkv21EO
zzgrICKIdg/EjCn2Rjp36gOXyms0+qonPQgN59tO2ptpl2DtuZ5ZCw1ENHhlVTvSWWQBlYl1p2O5
/C+o1IVhTtyxdS3/gXWAC2IVGDFUeFEK5cGzOix5XNRfjo1jBKsOnXNuo45fnmlt8IW7M0jOCYrO
wXGUyadt1Q/BKtZ45oiIdXhDG9B9NBuS9g0VRDo6KDfbUGTBUVGziotrV1tUDccKSs3zHXKYmFB9
OT9I3jPsPOcXpASFwC8GmF+RxT13VznfwmrJZO6gkmDqdIh77nbZdD4GROkVT11V7aJWYjYh3BW1
k7ofMuh9hpZg9SX8lw/NRF9fZ8jZtblNNhXfdAZBMOKEJYGSTdnr/eZDHAqqJkFNPRppkwuu4CFn
jg5hqAVRjb+z3MvPzZxcdChqAkWCUdxreyDjS8kkYTp7da8vnLm9H9SbX5LsnMKg+tGj21wsbYWi
EEvGLk3WWdkAe5aUQl7uFg6UtNRR2Q1UYnZdV34TkhNoL+9CWXpiCCATT/pmQHyog6jnLu5VquMP
afKa7Nmx+8+RW/iiyt1aKrIPAaSlphKkBC/lqXb8kaGDHUn2L+Jy73lI2wwU3dk9SmBTeBa49XTc
4RxiY8aPSB7ulZkmg+6Dft5d64eictzAoN9vy3fR/w09dLzMs6d2EpqNx6EYET4LXlOmx0L1N4nh
+5z85sRfTcTJBG+Jv7yZD0NwLQJF3VFxyaAGwpblLDAdk4wip3IhaE7jViHiKEzEFQAxW9x3r3dD
+0ahVeO2bjV1lG6EX+CB+vWb5W1cfg37QgH61uoLCI9SbbPL2dmU/BM05ZPaw6Pl+qaY73zcdfJc
1SS3tMfECcTzgDkdSh8LVWPlvyZWEnevDGEgEuRvt+1jkNcyv5G/pkeOHQ8PSXGqAEWQds3IX5f5
IilPnd6j708EFdcNS9yN9dhzlRJDM66UklZGOrBlUNuC555F00aHBXNHB3vpYYNx8J+Mv0y/DrCb
yZNdSky1hdat+9saGUkfGisTfgL4QPp4jslbMTDXMgyuf29z/zdPw3bjYRDMUORObUf4qUVr1k3C
BSQTuDthRsXBaonEeAh8c6RAbMMMBkFa0Btq39xhpEsJ3RBqVTNspWCjDpPDhy+9h73QnEV8381s
JxyPH8qWtiV7A95dCltvqYt0q1OaFssrCE5gDfRTPwkdAD/TNxQNU/Fey0rychkYiXTkFTQsDiht
iCa6ply4tGF1ODA/chUVKAE6ZA8gagbcwyvbigpviJSeBMUOWcmeBXRM3FKQXy2STX75YrDKl3Hq
kmWWqtb5TsH2M7Qp8PcW+01Sx07r5H7luwuNUbNI0KF+7VL7t3Bhp/30zb/n+CKCYevTSDYGCn3M
G+jC+8RAPGgReMRdZJLqXiLkn/7ub1xP1aPod6OFyjxJXLtj8ieajRttZ710rHELrKMCByX5qOGB
V/kXj9oIr6m4AxY6OV8cqzzEig6lXr6eC1zV64kp9Jji6dla9Q0ynPMuD2AU+NZaAFveCM4zv/pS
wTP2TAY6E47hVMxsLzFsJSUCfucMJ2hxXW8A8/DWWRzRu2ojFO5x0hBkOT+WQ21rU9jOX9BC7HiA
IzQDkKHdJzoUq1XgJoFGi8RqPOzTatvXx2ZEgFbyTcSssmwCRPgToqym/KFVbE9VvtEqIaMs1OB9
qdTOoX9TmrdyrbEAPNdZFQalJNVKHrCPFHuubloVKygrvWxaWmTvpde28HzS2s0NLCW+o295AYih
dOZOM+ru3ekD5N7UXKw4svWjLYkIzieDRV5WeMv7lN1R+i64wlSthS9glzi4WYeHec+tU9fqq8Sn
UIludEh9qV4pJY/u3gXAPhDpw1T88qxqEzUn/Jr4bR0xjm9hcTiIWVD8I1EgLIgIpZlFqcDGw5ZG
rqwjM7Suq/NnVgAS2MfeN6mCOzu+vDfnK0oKWlrpanrFRNRf3XbZVXkM79R/CWjt1f6LMBm9qKmx
0D/RlKVFDCqPrhGkNt7R6menUUvb+ferEjlM4d4i3NXC76qfRNslfykC4TdibkUvlfbRq4C4tUJB
7P3RiGGl6+tgG+z0CzNf/VS7nWsr42QteHHTU1T0Kjk0wpHpVUVFTUpVF2asN1soX87RzMf+Kk+U
g9EFrmYNSL4pjXHkLb7Z4O3iTAqu4CckCXD9JPU8ng67kigBBy2UVmRLRBcu6iSH+V/lJzmTKrRo
My0C+Alqy5uPUFUd9Id8BBEYIxsToHPlx72ihVnMTzuuc9Aewc+eetofaiGSRmHt8DORYQUjiI9O
29yJL3dWF/D8KfKpXMHcn6PUT5Rzc2wxn+TxJYPANnL5KVsWVkRUEpPoYElIMKUt7T9R6DX2FQCx
9d/1/u8kOc2A+1fPkW9IZkTl/iWT4SysFpYJMG/GzKhXEcKDIF9g8h1tl11ePLcDUD2DwJB5cLht
Vo/uABME2IVxoStgvDlEd1CCsUGZY+mw+SSNJ8CM+KihVQ16e17kLehYUYhkF+tKds2+N/ue8c9C
nVd5NH/Dtv8ovowelJf6tawZCNKAmRyrUo7u1lwpqmu/vxctAbQ2x286cJgjMxAw4yaoYggfUAx3
eUgCv7yzYS1VB7+4+C6ZU5tluMbreledgYH3oGP/0j5QKJmNzEZWJTo0x4JxHjwr9dJTtmDf9QZN
F96GWZK0212Oeo/9zGQI21aZp33jtGF09SSb2O64QdClxXSYbHJdKcc9WQhvaCb35MOK7VNbF6MC
Ck97+pWtrAA4mRjLFzkRBg+iGKkod5tkILaBw6kaK9ty5nErGKkPHUIfO9FUOXaL1Tb6RrUfEabY
fb7UVr1p7mg6uhkjLbJP71r1mfRec+jdRCnGXyay1XOSJ5+G46hiAy2mq4RxVzc/J8QhSbMf8AAg
BycqHvcGjnPwSa1PR61NooAM+iYtcxoYOoRMZiYSYhpbhbOLMqOnhWBpzaqLLCJhSOgP49ZOL/nB
ODorkI9Y8HfZWkOyM2shyRLH7w2gfXWXn4Bq1/ED/6kfHohlpVEqDRuRDfAG7J8kXKigHwVETR+Q
mc3uEdkau4VjwTqwwLb/HE6Vp9IcX8UUyyh++2C8cw/wyH8v7mz6/28l8Y5U3wBABjlhtBwkURkM
evsT31n+MNayxsv9FP80s8jaEZZlyo9oSmkdYcicu7Bj/MuMjtLiLsk0PXoe1CTZedZPj7nRxrHY
qbRcsK+e7BbtywUYVtPjGYFK2kauc4rIZ/lREFAHD+D6HsNgozNbIrY9GOAedw05hSXWU5xmQ+PK
Gy5xWCoyzKa23IRPvHZmyLlF9KNtm97iGJp8SBTjxTqhf++ydgLdmRKH2sURfKX7ha3zYI/yjpRM
K1KHnSn3cB4IpI0bHGawBSTWmK4lGFP9aBfEjC3nIqpN7BphtI8E0MGWeU4ZmDXNfJ+BWuG1Hctp
qJrMYL+X1FSGCoV2MnVS5XkS9Mtc0MJafZlnfhxPHOJvPEd9qqXR6V+GQ8OK/KaVbjvPmq+7Rpcg
ut5zhlaLsizVW1Sj4YcqsZuNnSR6j7BopOxG+r0OfAufnYL2NFJ2Gsf4gEmKKynozfiC2GW0JRdS
0h/8ouP1Omz1RYJqBEtrFIv9w2B0z2/IrXvW1ltbHfvNAOrSGAqhzgUBDLG8NZf2af9eYcDj/wnR
uQpBa84KbRyZNEaVGFqEq402/Kyu+/Z5SsGrbGZ+/dyIT9b69YYENA1Joqm/NT+a+bE54u1NjXr1
dommwNjJJPiZqpY5HHOJIdNpRMolu7fLpBQ+jbUhj6GvEpvwptnHtSeq7EogKCKCMMdvzIqh8uOt
Ia5RBXBg7iU2uPnGp8w755kSNTmwqObUiEdP+7QG6JMF4No8fTFuBEvfXB/f/xIntLZA7jhK6F7h
IyxbgP5WiWeLxQZ8sdzGtp9xIvO5Krj/H/kjZT7y2QYiUu/R88Hkbm7cpVgKcm37waopO/EzDAVP
ZI/l9JbKMSBiYcoHNiGD7+Y1kLMnJG5MTHTSDQH/jJnbwy5mn4g8BDOR95gWYAXLpBgXhi64K7GP
vLjBKScNnPADyiUPR8sZzS6REvKzEL5Z4S4I3NGh1hZU8RYlswFCFaRFvAP1VBDFWgy/DwOjh68w
j4qCQNqnAV6Nc5DI8byxWn2mJy/mnrhKDERF8MFLyIxfoPF0AEFhvSs/AfNFw5unwCLgu6h8H5Lp
Tulk3O3y09V8DG6sUD5aUNyT7Cs3/8R9EthXJn2snAkXDC/IodD2/iIZsSNbHrI5SqR9XUBm8txF
okAgZONLUkqHKJ8LtsCXpPRliZtudWJ9k82QIXnrlVkNX31oPZ5Yqktg5fLw9JXtzLHIkBozE3Fv
6wLm5heuvJiASULh5bpvVVUYI/Kp3BE2pgbzFL1ucUSX4ST/3m/g9QTWPJmh7uG8ez3iC4W3Ixm1
+vLjv93oM3kOz3lWxJe3ClXHLBRHy69r845Z3ybLcf44kW1nLYi4QyBKYDHlpDgZL0c/oEw4mqJ8
+TGmct5aalxR0bk0qeRhj42ZfUv444wMVm7TXnL3wuAAgMG4zMKZfIizZawCE7erDw6jRmsEINvv
D7dP08Jdt4fZ1MkK/W5M1gxkfMSINEWJ/Z1hvMLfGZJIqmKyMcxaTKkdQZpVyBUQjbCibdJ1IRtU
FITkrCa/kTuMA14LGBCtQ5rPyYgdsS2dBrdKO6vrMyisR9AdZJG6OgNFFH6RVGEghnn3pwtkvtbn
1dIZP7kaDoiDMXKbVWdOWwINlcbPnFvYr/0gXCcibtrlGRdFFyVaVk2WZwzpT1VFeXzY9aprpnwP
mueFZ4VRWBvPQzhtuvBbwO+oTpkXMjQsIrPqLfkF99E3f2NKk9MmRDLWthkV6lo6UynGd73ZXsxL
T5YGdWg5pSM6/VSKyCugF+f65YjXRNBXWg6lqp+Tw5hFsMZL7oILd7yvYOQK8zoSIG9QWG/ip2a3
c5hXL2aFp/3WkBSwEfy0hwBeZJW7eTEohA2KIFp8WcZIgUB3vSFaYkGQaKt7e8XnBtUch7vvCTrd
xKV2xMKBMrlc0akgx7kqEQY3lSuIBA4lWsBXrb4ruTG3nYx49Z/MqmVmGuk4Si+7Sh8h80wVTCDM
Cr+4VFPNmA780jC12oGHsnhJ9LJ2A6i8ktgbSixZHFwxODUasjwQrUWIwiETUsIsiWQ26WVaXYFR
x39AeBX0DMhb/E2m2EY5S2Qu7V2hLt9glH/iLbodewaP1YFnwBgbrH026wXKhi9GfxGNzS2Xpnmb
JEIvcmnv+SFbMtvzQhrVfzDplDWBJrC77qQiNj70P78BSvP8kM2UFQJigj8b5IFIPImvguhbMIms
lLSD1KHqd6/SnfKA9A8/S+zwMT0/Mzq3xytE/2wYbAetLIYviZesSTOUBrxCsnlV7Z4GMzeV5SjC
kOEMIrADubVjt2tdmmltWFN2L/Ow2KrGm+Fyphsqq1oWuC6vmxrA184gZzMZjApIBZBm9ZYW10k2
FMmqnxJkttFpHOeck38hPhgnXaH6DzNga8C7GzcKv3SuZOfb6OHKJi1CHqoIotbEzdG+NLOEgBc7
9X5YuMqrD71otV7XzHPhbgLhYhnxkg9rXmx2dUtljv253t/EWkwqAriCG8qC9z05QF7g16K25mZk
PetGsZlK1YNJKl08ctlmRH6gQ3CVIjrUSDpYEvXLr0n1uonOndxRqmRCq+8VIcwHCjEnwaD+/CWZ
D59JI3RaEfAUT3PEnPHPsIr0MYZYLUem8zq3LTprhZo2L7d54bpVklVxql6D+yr7tjGszFc0nDpY
mSVVXxlvm0BxgzbJwbP3kIPebgg8/fwNh9QULc4SXMae0frzjuAf5Wxt5yuQwRE4zCkjsXVKaJ8M
GuI6kuNvl7UYArH6kT0Dpr+kS/UWLRcigW1PJidJ+a3yD/LzlqomH+qDHlv5KKlaj5xbuk0oBk0A
pueB0xM5O7KfM0+BhV4mYgcQvbVhGxmnEmPSKQXpeZn7mqOc7tIN5Y/CtDa9hXqs4+5Z2NiGiYfA
HSulKed2PYwy0KpF9pAOyMvt6CBr8VKMNMor0bxX1vI0xxCTYEevAbtKZTDUgd5tG6jIOrKi6l4S
QJmIhk/QV4PmexhambfYMjbE6XLo7/9Eoz7Q53PyU75m62YlwSzctyJX3ye7vBG8V0I9FOLXntiC
xQ+IrLxlU+hnx4cPpGsMwzMeguVs+uTHaBxEdYf3PuBFQQCQl7o4eMOcVjFt8oImH1Lsl+IYlJPm
8mjhoZViFTt+ZDE9U0B/4lNelPDtmJFzu56hh7cDvZfJjxpRnDmhbuuoxIi+ELr04ZejaHUajW2U
SGGe1dYTz1zrjnxLPZ/thThGmAqfvO/qWPgDvP37BcEwI9O+coMk71as11brU4VHWwOnQeFVoTHX
9bcZFEUO3ODMFsnG9a9dS5TwyyVVusbVIbxFe/sMwfS3mhfurH/43EmeY/pcn8h2lv4LP1Uo6uB7
vrd/D9wxhcnj381OwpdRcVSozag9FBidHZpucHKHKchBeaHv3IdfC5pqqizbuSGcXHsUg1g/ruYi
Z1Me8fot0z391YYTjnr6a4kNOq5uQF6xgzTwTpln63CH5R6EXsaS7ZKZ137oeZ4XvjWqI+6NBQaa
4o8kwvnjIoa+rw9HoH5C0tVGefcFFiHXX4F+SC0kiYijO1ImKZF3qi1pDrNODIzoFQInhTmNAiVH
bEz6X9z867vZXF/LB1I3Scr0mj/xsvTEqrYPPP8yVGhDGt7DUKWkKRqCdcKo+eRGJGKe4CHB/0ZF
BGRGQtypgDS0FRNVJFB2NCL/sG72QBmAMEtQ0lKKTk0uGrVEZMeLUU/J97XJYoMBe3w5w4IwmdGC
sDecNKBbQXjNCxxXcInRQkEkCQ+YVazc4MdG05tz8F/cXlqmmF1vQTIx9fL0ygHr8KZ1XINABO9H
1pIUfXwJsmTTruX0wO0EQrRdq9artHxafC9jAikev9gVZaACAz7V2zkkWuK0DtjO5CiqJgDECO/j
YTJSjkGME/TP5c0IE4Mvbr9XIWqJVc1439ZIIKjmo8oRhyAvvsfMOI3rGgVJcLlE3KHPG5r9JIx/
PyHOVRNvT2DwqgzdQQU4/UhUTkwtj9tFqr+devrs9lSR2GHcxfhPgaVAQG31Pa7VQQzFtArF/LGb
2VZtTIWxLDKlYdNIHXWjXOYOer0aZaXLuz9Q32nY/oEpOfStx33Q02im2dHTYmRcI7XGEU0POXB0
PY2Wt1ML0vlKkeMlQkqpLk11fzgethC0pBQwPcyJwU5FEmIpBEkARLu/RSnj0BkxOlq7f4Wie5o5
tO0w7Ix+AMd5XDYj9LDaYPmdt8JT7aejP0/m1Z6+mIYBDzdC74rDR46NNrsf/64DHrFXrEQm8wib
VKYbnkNxQpNRSmVl4nUds2APKmydhJh1xXVUGGkyO7np4a5BArOaeL8ByyQD8A0nOMwxs88I4+4s
ovENQ9mkbtU9W/RuS3jVIxwHeqg4thWjmQcA5F6ZLFTdT9G4WD35wvTeFYO1EMz+aQhgFQD28rFc
hFdCuAft0keQmTpJs4NJJig2iDq2ucsyDd1yfhtZ4c9zkU2OtDcmdDt4vLb8s95Sc0juWX/OCRng
n+2dqG1N0nnnzWbbc4mGChyL/cgV7WC0IZEy3yyVjbkR9b2W8HPN4GilJdZtu2dQeoCk7ItyVfjd
G8awn6n8K5B9CHLRRSeTAvUMcVJ48lpApk8ZQ2+mF7nvUSpXyiYP0Gx2lbEruEnRpgEviaza8PLI
A5vfT7PCgNroeMLuxSQ1lpS0uwVq5lzgxh4lE+Hcun369Xz2T8SjK/E6q4Fef3bSadQLUhF1Ai8l
Hne3F4QDWK0ckyK0AXV9F0LMKR28gwKBP9c+hNTeum/o2t/SzALWrupSi9PoKnbKLOYCsVwUBED8
1EZgX6bkq77/hoMXhpjL7zzfIrseTdhoikvk8IyXs3VRNiobzcjK33eBONTc0mVA4FUkoiaTcSVj
U/XXfZk2P3V5xaMnzV4U7kuSyWXhR+FdTHufw9tpEAR7SVDNmp3Zi19KfehF714c8l2tSo//AJTe
cqcbIMBkwixw4aAJDXXKwYBwrFylefonlosMxVKHoIDm8v7u8XjbjlvJZBxESJcOHbemzr2cFFUd
E7A7gGpNtPUf62EzCluyx68ec7T47dRCxSMsuu/6lRKGRoULe3DBzyO+VKgIEpG2e8P4K/fnsqWQ
ILLz/ME2waAQ7EvIr8Zm46AT1eeca9gONldj+ENBvcmEV1WBg4tltRi7/1gPgKIQTgSaPObuyo+E
lkg9afHLA2o+Dn60MILyOsv2yOgl4voIpvxgPvzxepZH5t7E16B+6xS17/yEV9TlwF7SU3YCQ/Lb
TYns0rDFW0D+p5V818EfQZDHmbjnPpTVB4HZD28Evngo9rvDH8pP/fxgjimAlJAY1+oIz/u4biVh
GmVjgIk2CejVrwMFfVMhkgwbd21LlhM9aYHGAVUZbTEmz+PHriFCAtciTU9EB0UcjFFr3ZBcq6QW
PCHbzOHBbMzNHd4wqBe1/bWUwpLHubx/kbGkuqkR4sfZE1DHBMloYV8FdELEimLa1fzyCNA30ry/
z+hCZK2gpf54pHbwukNetvju+jCydQJXyxulIf5+3DAExzYJHgiLxK36hsGNIcX5Xlkpsgbu19++
HJ7qbPUXdg5BeXCnCXXq4Pi3p0HY+DqS10ot53uSC49ldNB+Z6WBIdJSHDzMFyWLw7bUAZ5BnfS/
tKdHECz2InbFB4HiNLvVfHVy5ue8hmEEYQFj3ngyLPEAKHgsbSYIZs1XDICK+r5mLz9cr7ql28s/
yL9a25iDbYN/Eduip73/HHhXJd0/ke57n+uWryMC/ZOcZUB98CGfNmybBI6j40vQNDrKyySEhGYW
OIffVaMmXZN1cFvrZ1LPCIU3gV9JauAm3PHJUfC3yrCVCg+/uueO5XY4pAc8r1ZrPbMCWqNQJ2Py
RJO79LrkW19AEir3ikOPqg2PYwVmQiBB+lvRXXSLX+erwdgam3KEIf0ZF6f2PI9kGhMnIzsh+wf5
ehkMs7Y17q+84rcaOyS1AEm7/aDnjubYCmuEI+7gFNBKoWiLEuh7+l2O9h3LM3UGUw03m3UDXT51
XEPir5sNZE7VXLnrn8Qq8c3YPnj6KwKH9rL9vxnxTmltbxWK0eIMxz6Z/kBv8q809wBCSeIDgh3T
GFW+hJfvfu2a1xnvGFHaCgeJN5yCX4FYwe/HWCtte14hwmWRYRMtQ7hR8a6ojydjr4v/yffBzVl/
UxE9u6d1NkOmqxu6ZCozbLKbJ49sMj6Zqk3su9HrrU1vmY+yZ2mao47/+cek2yx7cB2RbauPYfdh
98xLZnjeDIOsreKwCqrEje8tBAAAB+GILRe+7LwsKIBYZBzmkhv3UmDfX8LRCmylidKYv1D6QlfX
ct6E/1/NLFcbVITkdElmoUxDImUptskXFPGS8FtpTDhg1r20X8AoTdE86E49O3sAROy+IsIVIGYz
NzMI6727emzQca0kUHe99BUmTSb7qcWBa7CyD6jwp6oxwgM+LJiQw21t5m17E9jGMIvwHFKO6lWl
FCGlU2CdnWk8dosF/Jz5qEgMlJHo2FgJx4bgchkxogBQ+U8pXYJV5N85sfBvdrhTZTNBCUujxuCe
WB5ODQNm1RK2TwtBNvtGS3kqIE+IF+P1fYxcToI9Zm5jtHQcC2CSMn+8x1vxyRkygwPjmcs+xOBr
tWIkMaehRe8W0QGPhzAyYcVhmZi/LTm34KNkYofJ6U3NZMAKSG4BCXfsjBbj3tcQ0wYwM/mtULOD
G0whRjK1T3zi8RGe3Tew77JlLS+BWH5gAyHxB1YBZu+xJzQLIT1a5HGLMdSAEMvwrlAfK2NMkcnM
7CBn+iKmPLBYofAhPgqyFY9jd/Jo03WZPEHjDyTJF06pdJOprWswtB4JvKU2Tm0cNFnqnSBUZaE7
xIW3IOsdaq59p5GDbzG5weAfU9vxIfEEiZ+dlCnf2yF90pwneKUI7ZFLf6MBanCe6b/oXZ4Wywse
c6t+d+5mIda/9I/9vXj92y5j7kD1JReKG9kOBYXhlBuhVl/CPle7XsInOpbXoHlkc0c3VgpKltCx
AxTmJFH6JAOA8Gp+2XY6DAN5C4QYucusU5wmZ7PM0n4NELqEeFhC8s45Ri7wiczWJ1+pjz7zO3WG
7hpDC/tsbgxeV4YBS2vwmU4JnerHwdq608C0inPg2WhPaYh8/HVuNpVxd/NF3qcEPyrqVCska3mm
DXyrpUY+oERSIZTehclfTdl4haUB3336qnT5ECyAxiEXA7jNyNTR/Rv+ohlToGcQ4m95BRLCIAbn
23Uepy5kzn6Tvaw7UxFIaoSvvQNbh57QqjPxKR39Ybob7zuQfxdaREL/veJMrNIMW8K/uPB0umpH
ZQRpZDKn/ye6m2D/GePn4/sQUyCllizKZKSKR4oRjKqYdiFssgMfuN+iCB0Jsw35yALuXvAQyiF1
R7xzq4cBlfH78+I6q7izeiN0rMUYTT9rjJ+q+6aux6ORlUXzsjyWUxgU3/L8cSGXmNWeROAxvITF
WTnC8puGJNjNHhSgqkBHSk20HL1O3nyobKCfEesgBtUHUqHt+5ZuS9gDgYvaNUmuNAQEv9CF/Wnl
/GCudxPwoJ+HrGNfUfT/MRqZQ7T4J/j/1n8nYoCWM8oC5GWFLN2DR4FVz68FGNoJRkH4IRav9SuE
ME9Gm+sYkcf/XWquQ22c0joJnk8pm3OM90cvE8klJmtO6pd65A2WI4SpriX63cEdy/aztoaIA79b
4hH/IeG5Qc6aBtmOQfjLN7sTwCL5t0+fYooStoQ0+jr4HeGOzIW9MGFGOWEp2P9o/qQQUoi9XxyT
+kLTPHn6yz6cwWn3OVkFHlzciL33OvApW9FUP6x2P0jbiryilcsjiDioaL3ta/j+3rbhwle0JH//
4k49Igtb/Mnr2P9AOnJOaJ85PDVL666gHh2NDKDehBt0KX9PfRl8KyC7WHbrSmmAYcZ6dlsxYyWc
Yet8WBjqP10wju0P7wAlV8XzfoAvVhiF3T5UO553i7SoSBtnqMXmWki8YIckXLuaixnxzlte3Ddk
LZjEZ3isUdpaoBccJKnl2dZ2Ii7sZ6+vzORDL0HPaQYYkSRq97N/a99XJCpvfTE2GHxxbT7V52+T
vTK4pd/N0ssDtc0tfop+MfLizZAL4CrjS04berCBZtnGIMMOGcuto+oioF/66oNT2/9v5w41BFrs
3O6dJfDR/tq/jHRHtLFRgG/l61Z3HxBNNSfY6rKjnFa6Gk7btY4MvfgstH2IrfkBpPuL0RGkhtJs
UpNzkeBbON22YOEPJ3K9bIQ9K/aQn+cIUnnUnjVFZ1ylbpNSBSivHUiquuDMsfPix92YHsraHfMk
G1ICsvsb38geOxIHTyVzw10UvgtF/fw+eZwkIeIIyiQdy0/DVQjRU0Omhntawl8YATVZwlSjmh46
RNGLYUANKNDx6FjgA3XNs68ni30k7lJwDPRmRHpoDEfbX2LMfDfWvHMgQTHZ8MtBOsOozhqWb/a6
DeTKgjTzSmmdY9JhH2uIgtb+3FrYj9vo5qbtdA3tC9r4LBRYLnSrjmXLfvyoPLdhugP4ZVcuHQDF
n0dHbvJTswAz7uIzK1paT2y3bF4/8R7gx+zv1u4FFvQ47Ekpsg4hiO044a2+oVCyYJtecE4P2App
1KnsmUpvJ1Xsuk4Fz8AVk1+84sgJ/FK6Jn+VVtWBI0Kttw3vUsjw+fYVYU87T1tPHmzMS9SbssXg
7JZqW8Tg6oXUOMpHB0XiutwUUpL2NAj3sK5f9jPp7s73deOPXXgoX7G1ckqTW7aepOYid4CXnsLo
7YbIKIYlypXB1k0Hco4Ty02lkEEN1crAh+0g/7DbcaPRjm0Mj9LeZjzXeWsqfTz9MrNU8/iTBIK/
kscRDQgSDkkWIbtIApLeKc2xsosxwZGuhlFGIRkLb1QRkYBdRVP6ORwxc3pIDbFLnCpIVEh19gKc
rknFcQ45BE1fxYFgK2quCYKgeFlSVf7w92tWbEaliQWbKHaR3+BVfb4zTiD4xHsF4z9RQcjpS5Z7
E5ylU4j87uJ8/XqpP6NEQ/Iu7rOfHCiEtHfVYULd1A3VsauudcOU07ZBJzdGKWXrNhjdo1XdGr5Q
haTR49v5qyBAv2doYBMl+CcoOzGPVjnJLmM90wLW8EuvRv5AYfdH1zMPQLRjHiFYh7Jvdu3OZOs6
pR7qHkLw3qfdiXh0pFi8rGTAIPP/6jtgEIBH8BMyHv5jcVlNEHV7VX/7NAGFQcJ7H372rhVLn5gs
TJYdS4J4+a45Qg6qkeexWrVxkENJ7W4/zfxJAQS5mhonixvBfERLQtWF/Nj6TJUF1cgEb8M8DaOe
aY6rf7mMtwgBBSQ9rx6ik/dRXTlEWGlEgRSfDbILzhrJugvBbpGEmR3rspuAsa2v0fVh+XGKozwv
H0FQjhpRbdzux2m/EN94meQvXYyEQxERKp3dp7irGyneQcV5RbL+IV2ucu8icHgG0u5C+QitvDeU
fQZVioDwZYl+EV3X6WVDJdqv+t2meWbis+4/GK157vbQ9j2TLceK4HhqTIfYC086WBQSVjw+E6Er
MLy0xGrpMc2IvBWwTdiakt4Bben7psdYWFBlsSVgw/64PR88KAq8LtpYyKq0Uz3FVgMhoH57n0tm
Kfs1VxSLRdJKLaFx7VdiI1O5JaCp3p1RTHA1EKua2lSbPPU9+aHIUNTegDocnqR+wpeBvTrsS9jE
+mDnkNQ8YDCzqVaMMEhlcMKL8UUpXOQu/rfG7TyeFQNggmExfmuH1K72yl+xJ8PGfb/Gr1hiNlbj
3by0nucFBaW+q9+0XkagP+ZGj9tKTLPiCZJ/UMFHTRBBvudoL0QFm5JlercAi7sDwmr29FMFVtI6
4vQXVbdCmg1KVrZp8ZOSvjeTict3APFMVMJXZ5zwMcbkH5O6NV2uuHjKGFoBhIWqWhmyHRn58+zo
lt4+KYvk+RLXcwnI3B8FPb8WWWU9COMaHhGJhBI5bxDudtUndmua4Gs+LJjYhycttawCf29A8JRk
3JHHZN0qFeU2TgTuU1CCJmJfSsLlfuAMCM7RjmcS/HsBtRuw1+RY7n66aZZR7fGr2rdQ8SaKmrUc
V5VsVxzGBgi/JIJTwEyrw5bDUI8C7lHoAt2dYSkpkYnpQnpST0TpHIARXKzp6EjmB7gLHf1LJ+LB
LYTC54Dja/nZuDclkjyuoFJURheF3YZ6QQ4dIVKifZ1T9YfEytsGBitLQKTl3hFIgq+ZyMUnZ2Ll
yct0Vopo1q25FvEsnNketx2HNu4TDbTYsa8HbCsQkKci8WFqSfq1XORpxy/W/U0gVQh/I/ZulXLI
bF6bAsSMabXloBEgABle0UCw2iRsrvFd+/xuXlzZ1y6WAknFKIKR4BxzYPZJi8HG+UFX5MCBk3WN
1yZZsyryRAzftOxh6gdB2ATZwteXdt4ydKE30iXpHDtYW0cJe4Pu8O48NC+r4OJ+QTl6ASz6gio3
4gd08TkOYpzQyDxwOKeQHUQPYTe80ILTqeTw5bjdWEq4lRgzrl/cD/n/vQA03orOSgPiUcp2zNdH
gQeBeMtmE5NFrYniu00uyBL571b3J9aG8snEYcjK4OEuAmvINbenjxybG62ekcMtEtTbav5x79dX
QRtKJXlbKZw7OM0yGUlQSMs17eA5BMTBZn5C381bZn0+TalZKdwUOUSFfAExh3sLcdK+x4M1OYQi
Uzea4bPpe/GahxeD5/PVqLdCJIf7buMdLKPJkyC06+hoz1TRyhJYqEQMRrEfwj/CDC2/1ZCz0JLU
mCcU8/lXbziS879XZd9LFICZORLaWSmsiBvsK9bpp5DmPrBenhl/A6PkyiWdAUx1HxGHl6DK+LC/
6swN0m6tgqyFs6orgaoH/YTGe1d3EaqY19UBfPFWzzy7vE2NI2KUBtaKn9xmRxYdGoN6kPF9GPPm
JmRyiSTE+aOtARL0Tuq7ru0E3iaSIZWzyN6RwsFREMlsDtlhC3qYGxgLnlpVjyYW4QqOHH7ppJmT
UR3m2FKJikS5xHmsHRauqwg1u4zPIcYUUJ0Z5gQFVI5w6i3vxEke4ZsRLKHLYaigyUyFNjmLz+mI
J6rbDFEbxuQ4ZMhCzNi42jepEad0D2rwys4ebo89Pw5THyXqMw2KbRTZm1tO9SnzbmuHaX7FynLK
Xd8p7MCGUzjpp2kBAR0ufTn8+nDeo/urcMoHOEpbBw7YMDhGCqSLUbAtHakCyGMAejg72yVasbIu
zFoeOs1AXZ6wmQLJW+ExIcyWi1VXq34VB5A917gypE9ermgwmBClJ+kvOA1EkL2AIXF+/GREppov
rca5+8wBS/mSs9883uGuukP1piW2kAAMh3WZC+WI3DbVT7JAbBV6h2uDyKFTeOmlH4IbjBsC6fF7
sNz1N8ofODjtqflBDkByEYnp0LFPF8IAImnWP+hUTzvoXnThqcmqHsxAh8Kf5XUIEtolosryhaa6
LGf/PuvU0v4N6he+BN8MjEF/rjiYYK1QJ3AT6SgcQ/u7W5VML4Jh30ctNrELah28gviP7olv05Rp
3NZy/rBod+WUJI7HlGStXUexa+6bZtOC1FcLiG8tF6HFoH0lz/7sm3+VesakG36lDgdhHVygwWfb
23mw3thhi2rnoh6D+lVGNA7U5j84vA0OjvNKVK4WUMuHW4Y8v3x/ekqkUhj0JcZw8EbBaa+PJWvH
pbHxpnPTtheQi5Vn2g7wFqHks/uCPQb7wfM1LmQnfML1x9uNulNCrfkBWUDka06eUtMTTvzIGdm1
yLBOrZxBj3tQNE7uk7YlKLzBgidGKwIY6QdI2RYB+SCqH85edZKR2fSkvv0avJve/XdyuRJpqeUY
SvvlAzPYAOEC+YAiaiZKqFZaqZrhAnQo3Monawx7xDai0RjNL0ZpVYNJFOMeFu250q32XVD8DF3U
1qgHlW2+2RTHnhqloxGgjW2+YmvAmw9XuiueXqih1LpS7ANlA5w4XeT/yXz9sajKm/ZwOAUQJJmA
TDmAjwWjUkA6u3qBTu6aH6PO74C6v8qBWaUg8TESvLMLzZ5xD+qXdq2TKqX1WzqTYhXHZzwwsjnY
r9JFmC/Tug4VNI7jazobBSL87k/w8r2tyRfjogazZSrQcmwAYcar/h3GaqaUQxXIG/L5Cd43rsaD
d48u5LtR9hVmkI8uKc5HTQtH3gIHZ0ED+QIdi4U+3wfd6ZEZqvPmWt1ESVwWdaVX8xOa1qlLtg7x
DYnhJwc7GJxo3bp3GfGrWSJbPf5mxuLsG1pED9i7N/R43f3ExLR4B3FIZd35tDHSp5Zb+fvIOUD6
QKc9SpUjmKKyaB0f/skjFsaWcSYT0Ad1un80dRYScVRs5eeT5Fa/fmIcKJbXcErA05+Kkf5/Dp+0
988UpxfsTEMYcNrk/0hL+JI94x7U2ZkV+VsTXzZ5JJMeDgUdklHg3Tw/1RO9xUHgUfVhV+RIBMiY
VjFTJVRW4xU3OMLMjqfo42GfCKJM/HGHy1kCec2SLfk8TOWrhgeXSEtU6rM95eRwoQ2OTsuegQ2Y
OGhFQu3pD7fflni/FV2V6RcaVMt+o8Hdfvv2HlQzoaqbtSyQGmveYcHK9vfTEmCx7a/eMboHDgZX
c0Tn1aGYExq8Lru5pEl9ihmHZJrgT4qORUdZ9lb41bEKpwxsd/gljUnlw54+jy38r+aepKFG26JM
ZGzt4zpYigg9WKxWQeDfKd+OESgy8PBa6HL77ofxwf0mU2W8Vct4xoEj6QPapUG0sK0BLOxk7RXG
EsNYxXV1zvZBcCDeTUU8C+3H7pd6h3l7A8SvsGwrOKKKft+oN+OEDYV3MJlRW2Wd/MQrMnmH61BS
axzyvNqHi58ZIoA13tRTu+6mJqcyeMHrVTvq2Pmfh0j28yp8zBv6OGsT3zST54RZWFN/1Ai+/Cc5
gcVVSSAh7iY0zIQ/E/nTqxFgq7BWYm2cl5h/T+Sq5zTDB7sc5Wge0Y8u7fC6UtpnoCAWJ/jx8awJ
NxPMct/zDePOz6f3WR450c3LyY+pl7XJpEZgMstyW9Jxj/xYE7rBC/0RRzAUk6lJAQiZbSdIYY6L
mUMAayDRHqyKPnL+KcOznx5vM5jUwT6qfKyyA2t5uczDvBBQ5fRrN2rUYmjqCazr+P7paJiDDRfh
fENsddUpBI13/ykDlbtsgO+PWaIuF2nWs4+v+u6xydnxQ5XAT/fGV32b1Ji24srIpLIV7MdLz5H/
hDX4U0xRORYsjQ2TYwQ68a4pSeb1zfqGuwIa9Mt5lhqXYqpyPeIotl1gASBl4Fm/jdCrP0UwYtUl
KOVtjQHPzkoyEqiSZxoccu/g0J0OZ4dR2urizu6T8sLxyIjajbXFMgViAFvF6xQWgbFG8gW+HkcI
ZkmB21un9A0iS076KfGiUlLBA4e+89WOII5gT29D3Lu5mvB9H/du8BIdTdimT0nAoWC5HG1TPDsa
MmrvO7teOEAlqRzuRPm/ILcTWznLl7Lzmap5C1NyuX7aQyS/l+Us2JlzCZmPLE7yr/OpE0kfT/lR
bAQqkuZAhtDqhwmCtZYvnNY3ipZkaeuc0hjg6xLo6DOCGwI/qRowvTPLrMiXBRKuLsO9cXtGI7Mn
NdhJNntDCbT17J1L8fFwOHZkEllRZJeVCOlcEglZgeQknskcTAvYviVfM8OHVfpuyMsOc1oGaYn5
i0AxtRsuGGv7K7mcjZoCB8IkUpyv+ksBDAehyVEEH68Zg6UUIn8atLIjxKr2FMDJwrWFQHksVCvk
a0wTH6oWemk+yTNX1T9oXw6+//E0k2AHo8NBGwqtgcGOJnRGrs4VEnlZby3MhUeeBOL2jU7CGLhw
o9Yq1/EeQHgOTOYKs84QTueFjhJsqGtxHqvMt9lk6zCc01XIRvtOhrEOHhND5tTTKYj+RF9x2D78
u9Oq403k02sVkjrRzn0z19D0qvc4faP2DyPtWXjCrpaS6Es5KBPB9SZfvpyClJ/2vod0Utm6Ce2V
7zPC9L36c1t+czqc3/GW3JT9dIdA/vQIMflL58ZDV8E3SCdBIn1zeivYV6Lxc69vrMHbTwlypGIK
ovVVyA+XEwOpjEGUkhA1w8+dhTK4qNQ6h4tV/6WgccveoqOtaTWkrAMj3eZsyIm0aUWj1wlF2Bhd
whXML3ucC5CsqrR6pQ5R6dnfUFCjANfLB4V0XbgjaPsQhz7x/w61Rn4noQcyNOHVto4mg4Rt9ad+
pS6G0qBk2bWPFq4BNOpLn7bwkecH8m+xCFQiGSE4itBdMYVfcY/C2iWIhohPTYNxvos49XFNhw2K
Q1jAEsj8tTptwAlyvpSZAXAgYohMU0huRRK9kYMpaP/yBAfAA05Ayo5FFU+xwhR1yQSbi3rSz+M/
gqO/XJ4QT0um7R/O9RdS8kH9ctlSl/dy99AMdjFhIpLLN3Omiu9b4UV6uWWRREG9QMdiJxQUVaQF
JGhSy6s4y5+Rzn0OSQopztJ38MlJmxkRXvYgqKpnLFXL6rLLjEGziaTQTexBcts2OFCd9eTT4Sab
cwPjJLBzc4cmoVssE+aeI+yW/buKxeAkqXUAAS4ZQsxo0bbaHsP+JQFbsJ6xDV6umBhoC4KlPNTr
p1yz6hw9KjP7qhT9lytmmm11Ly1ia5c9W47GUoBpv7tJCsu9mCZB8GEnxRR6wHgj7ieMY1oBy4KJ
wTGz+xSpBVum5OHlVDhOXvvk041YP1fV3UohVpFTREbUvVdo1YKBSEGiNK8OgrmRaomhPkBdfUcm
LlYo4RtFWsxlrhanyhNV01VuitYITR95F9QBE38NUGg7D4wJ4TuzgjkQotqSkMCUVHl+o6SOyJU3
3jPDAHlCcIeqNqXjHZqlY+XVOailqLL704brI4iuI0cGUlnZLr/8ZfYxTm7p1yNdbODSd7krWCWp
vgtMztK5thlq05X50xfsx7Z0yDA9Q3+3LhFncefRo5TgKWSqQ3jSoPloRZMQpu0MkHYDgikpW3+7
cpB6Mn4iH7vF4Y9SHrBRxdcyHdvOSBO26/DpYJUu1d75hM4f0nt7agCo8A5odLYjHjAqkvldtkfz
Ah1H8LS0s/d2ak3k0v8G+YpVFpJYM1z7wUgbHB1g54iAajBmPGQpFj4OEHbfslH1wbKwOG4u128I
lYp+ClyUXzQhmZczhWUDnUo8pcg1OSY2EgaxdheNPHc27Wj0a+k6GRVp15HMVeCpsLWHwv3z7DjR
0Jg4SY8xVLOJ0QUQvd1P3KJzyFwlKyvzoSSmyJsSs0/T1pQqUDFrown5hMcZ6dHqs9YGgrIJo2RE
CynkeTZp0KLKi6K0UONRWKreISOQgmT5VfFqLzZWuIztVdhlpKcu7sNAdXMtJfG6MWNoTi5Rj1eu
QH6W3NbreW1Uqk9M99Tua+KLR/1g+j4OMgoWy21dGpj7DZahwDveEvfS6iFKZNP1PT+PEkrerYLt
6Mg8HcxOppiIPFxpU1QZAqeFpKaEQv9sFc9P2bBRV7pL4AfXGXKLNl05Dj/2+IBrgC0PoJ2PJu0U
LEthApShhlSMMkcEpaMYy+eYz1+tVQkk5BGXWPYPzoniIs9pxX3Kxznirci65LH0dq7hr+biDZH+
GtCXx9cucTXEQVh+Qo4mxEYCnN2f+2we4uxPxxRHDozvmlXbfgURK8hBRa68ySq1yReJEfyhrud4
lmnl5lRTNa/UDG84Ng+1SH780PQDMYlagUcHDcIkBsOWfqKytmHxKumauJqfvnuG5BymDGeBeQUg
ZnQ5u1SiF4Ld8JFsxm4NzyATUh9xGBNu0oRbjxTww9RfzQ1p4dk4vKKrXUWdH9+nnbVrTiZOuGMI
6tonYlZ2/kKJGbT5mRQtccxuCKMoDBY2g6bjRUxCuWZ0zetilY13T7H+Vc8VrrNa+pA7ULASNrL7
qkondSkIFXqm+0JoEGAC50NKmUMUpHenfkJ/BPVAikO63XGISzxMCjXmcqtUQ5aEvahsTfoo7UTu
xdtqidnbpagBQky70yqCMGv1lGfUXLMWjZ+2Z8JkfiKnhP4YWaARTjqysAQDUZYOLYoqqakFR6AA
ryxm63AAfGg33Cdwf9neiLIrpAsmmxSOaUJkQub9dTRQTFhKgdMPu601HSYDAHMznrQ0+GPTKLEm
RHjROW5lwNoTZLBb4rA5Q8MkpUXU2l+Re2Ac2EjTUMFCCqAnqeshbQVgsBSSZso8uXY4LxktW/85
H6QtYA8YlrYLieCRJ7U4A3s4bl2JtIyPqSqj0IupQwZCkfUNuQNAtEjbNUv5RLzEz0ZRb/thcKEF
f2XIo2TjtIuedb79qaeGBAB3hXQQx4VnWAZK8fu50F5neFgx8jN3nyGqXcG/IUuamc+CD7c3DaAa
EDrwHpMkFDSr9vDsbM9IhLDr0to8IPPb0zn6WO2A1G2KaRsXv2H8XKh5uGBNxiUMG62okcDs8xXM
53oTfPYUAMePykbJsoXWQerkjohGfPfTlsJJ6w9ToKRBwwXSUUIh0golj+ggWgZ+09Hkx9tYuomy
b+Sqi0Kkdygnmi7rxJvUPPv2UGNaoK4DzySzRvsp6Rv3NioI3FoUnHqZxpv8XMElTILn/cdLxhce
RbuxB7Gm1IO/2YAVsi/acPxshpcGAG9loHBDVbswnEiuJEES/vya9xeuemCZpnrk7w6qxvxUNLKK
h/Gt8fe2RFFV9rmaJ+dwngI0/tFopBW1fhQ6akDX8d+WRme8FPTj4qghjf2fbosKTDIcuZivE3GQ
AZ8okNigukvmacYKo/JxV7ynJYCvOU16twM9g8nsx9sgP9FwNXujDwRIwXIZ13j8BEGVf1SEqfQA
dEesBUmmpS2C15/KLxTDnX7DCE0LapSK08af+UZE+jMoAnWA68OI87fxRK528UFIu09HrKEWJ1/e
A8f1ut84Zf31pAlY+eWnMCddc0foOS42SA2xo1wLmpBs0Z39Hjkhf9e1GDTPR++DkVnj799gayE6
053ifBcaVITETBB2sDbnOmQ9F+y8ieNlJffqt2TUp1TTgUhqJ7uDod1qFt8VnMs6iez0TwC0cZqH
o0/n8Ed4tLXft8SS/o6d30U5YqTJ3sJXO0XdYOlKsvqpc3VFzbHvakUuk9nxiSJQJnRBF9GhcLjO
FVBIMU2YbgbnWxyum2FykNrAPDNihHfr6QAyE57ZzhWmfb1+nt9Gyczn6O27Kp3i2Zz8F10oxEMW
roquLTdR+7HiSetUnQXt016qcUIpGihCkowjLkeus/QG+MHAF6Q48u5rnGpvJNnTSx8kfIDoA6Em
QxOyQ1NQgt6JKW17/4ZNonr6LyXbbtg7LhZbzum280XnWOqO2r65jKe6Ht4QQCJOJuUPI0kRowj8
MNM9J8QWn/+vQlT2jkJzpJaLij/6PUxnGz4+vIgXRLc04c6qgq5JoBqx83yDaqlU+BjivmPz9mGT
cFKso1AqJxDFcTEzkGdQuweRSnf8r3ABfRW/YusXoKb9TMEHw55Kql08fAguhxnFC9m7JFI7n+bV
r5SI+MgUUuoeokv79LWg99aSniYdWv4nfOxh3EDjKHJs+iz8Nfs83fCVsgE7mRTRXK55Zo0lHGA9
8PK8+m6PNNJpdzmqcQI+bfFYMF5g4+DhGOxP8U2zG1Vbcl5DCJhJ5WhnFMV3Bp9VJuESMjxPkLOn
6ZuYoCUNByqBBp+60IBAijvGh65a0GwXTufLqjyGrn+2kaJyM6PESJf2/SyrIiTCGICFprP7XQaJ
lBx+3XhgvT7oX46t9ClJMflD4kYlD2rGEMq2H4MZnGXzr54S1WGE9Q1rfwz7WYx71wSJKH4/Ux82
Rsfd/EFI5+FOzD78WOUoLB5N7JJJkeRzfNscwVsxHhmDieykwC3L80xHNXMHrWuhpl8zHZVy3VHG
7qb5y3OEMiRPXnUwTrcgJkr+Nhe9pMj41LNP2FB5VlGpTPOrY0nC8X5qNuxiGD/Ce87RcSs2EFXe
sCJ6DEqFAPmxhVevbvRP88owDA0+A4u3Bze2lwRA2EeXYWozONYkk5oDwvOk2h6i80nAwLFquwXB
ChLJ6TjjHHfOJQgcptz7SaDB0+ZvOp340QA8YSe4VVVHvRm2LMZWKzRruzdz/OnvvB4xmmVB/kqm
lw1Y+zUSkET/wFFevV9aGZ517A81BNJZAbB1dryEzC0cOLlcoNrkwBvPOWUUeDD3x5Dg/bGQ3t7r
hMauSPcMOczvOyQGQrIsCJWUWO6loNdVXkuIL/sbfeXqnCm2VS40n1B+7oUFywk3tRIDE1icdZeZ
gyi+6RxtaJxolm31Blr6MbbfkQ9fmNdVB9091xi0l4O1vb3sZnonXHgf/OStbY51eP3lo4poEB8q
8VMLr6K8KRozudhKaa6a0HjMK/LXReYl61logfHGeyFGeeqMqjVqX30MCYUFv/aIhp9+8DjhA7r5
YrQujD5AJtt0xgZk5fYoPmXwOhaNJul82U5mK9q3TDeaqmRrAcrkGEoh4/CRT9vAcQaxh8fXf9ti
4FD7lCHcfAO2jx9kPGJYQSTqokEYyQMLv7/UMLdnWup0Tt7Nrl/fpN2WzB99rzBoKRgs1GZug9IZ
/IZTs/gpT3iv8ZKK5o/6nSFuVS4H3+0f0fDceFssrzGeBI/tVANuuEpCeXtFHAeAtvdV97hfspBM
xpaAgTr/YjpLIOuZIZAAPqLSmsrrPApJ28H15evS37WfR7xHPpDzwrsT/TkChFpXWAywNto8ahgf
+URg8+mRXfBGDTtKeTkrVU93vEtTqxA9XwC+ek+guiuZEQYVPV1VEbpoTYbvbaG4RIfypTX8YKL9
K5g1Vltr8QCClvJMtUCJPEo5ITQ/0eAjwcNhqxFOVTh5Ve9wpt0Ant7jWaTAUuJRz/bBNZXx8mz1
jjDv/+4z1nSy/2gJeDYk3pqHqT1PN8gJ5BULSiGLapeDRiJt7Hdzo/6/fn9zeGVISZ2xqY3Ywfym
J3yRvTWWK+KqEtdv4vYz0G0r5WqDh5+bI5g/wI87DIMGi+GUuH1AIjZD9x+/djrSCTFldpTnG2Qi
PB6hMwJ/mcDmLLlIHKCxNePD5z9lX98M0BO91hMBB0jo56LrpOe2uvEeOjW8xD0LCxutbp98TWq+
DfeYIKrcKf7mpTKQzdwCiuPMLxzkGrk/+RyrRIZ3fttvH8JEerO9fzcQoerQpMGeWqsN5K4YME0Y
i0Kjuc06A2yaDhB9gD9vAiFYOyl19M0G7RZAIrZQT2Ve7fjZVOpX1B5H4diyaCKc/4/l5AFF0H+N
/2nnU16wDNU7J0jm02kJ4SAKSJ8lMl7Zz2m8OZf9dHJhNo4NkGZQ7WgsO9VXHVntlOT/1u0QmBf2
ifaM342YbYJebDNWSD1DfuiseDSxDzQN//uYGR7bfuhSbbMHbH3CgMkxj0PmYy2tm9p++Aq2uZI6
cZT8TvHtygffHe5Xb0yeySejwHp1vp+xaC0EnN7h4kW9OnV6JOcyfsHAqb9g2yvCKq+NWFy1TvqG
cxGWZtaTaxkvelSL2MCUEvUNt6FliHMKDR3UAeLPb9734LUsF1yVCh/iJ3SS6ihgzWKX5eOcIdnj
mUSuAMkdb2KYodyF5Df6sguLWtTNNalgct53nDvvBOT+BKaM/slwquvOPqPC7wRN0rmve4XYcbTX
HGrTVtDLFMBBIVAERgSxaZgzmAi4TV+/nxnuV8E7M0CDmugb8rptY/KKBLEFGsbuhGPubhVAF8zr
YYffpTJSU4VneUxEIUV14Fh8eRjWb+/hvTWoRHn8Z2OXnIRdBkP93/0HwvmXR9uGhXdqxedz6bX1
jtBHTvP08orcpdHGVaLGb5e7HcfOykVcNgr7pyuZTyGMkWUSDj3ZcT99YvOBvs/12fjgNfYr4Tcr
95fpKvb7KLiwFoXq8TeAVQ2h71t2GPMypNvuxpKRc8uY/15uyNkN8QOnrGGHns/u35tJXICjacDP
ZGfj6j7NCGXvrKKikI9LVqi6/kXKToPwPCapbNoZe2/YOvOAm3mf5BKrRUf9CMRjRmEukD2/12N1
ZiDvAWZ02eq+oE0WnLjdiI8CzoylWBJYbx5ag3Efgu+RrMpobtwC7k3HLPAYGQBiv8p1EJSOJ75G
XG76Mx26gihvaBkCOyhWi9i/+JDungzK8Qi5NxJmTBtT60JGSCiCr+wPzm3Ih5Ur2YFY02DKUPSH
uXd35V/1nBF1byXFFJJzDYQjMlgBLv2M6AOizhLbKWmPpjTk616+wupdoV1OPLwAY1IXsZxYxFAV
v9eSod+GUXMWR7T36MECOgPe41W2qm1fQt4LflagixFyWXmhuW5XT/CdKpBSEMKOQYCqiNJBFiQp
uZyMhAFSDokVSnz0Sm8vY1mlLe1FbcoVyrnEElkP5vSqZNGjYpxGAK+DmMuDxOMyK1deqnOMlvVG
GgqG0aVryyVYXC+apvp9+fhZolxxFwt1R8KaL/KnXtfCGHUE0aGZ5uHY96snjV2oQGQTaIphXyC4
y1ixADx5eryjmjJ+i4eSJAt7xBqg83AjAT0dHDh2oowWChARoKRZe8RMHfConsxM1Lm5/jeMzyms
873Jk892TbX2tpwVPJwIKKBzmomfLhpZW6+rp+4mpdAh/LDSrI9yoNYCOF1mN2GnBhLy+A5d+5kT
TgRQRjnqOr8YCzd5UQ6GJlNG+rSCwXasf7KZDa/I5S7qhm2BmRCgPNkFUN4giCx58QAdZFZzFvpl
l9QhR2mYA2cJw7Q7S/aJfF7Obdk/RpjtwvZVWxGl0NYk2Jp5jiY35fUjuYBOpCMjqNUUunIm2uWq
Q5ifNaqs//JURuFibg0jFCGVQegHICpzxP8U5KFaKQm0L/Pe8qXYN53kuTkIyUnhcP3brgAv4q0p
IwWeAohsA9uCB5dgPPuWOQVK7ZRakLCHq9DQNP+szGx94N+uJtvYyHwDZ6Vbz0RFAGzZ2F1NzA3W
OcMzhkCIKY2jvM0jZRK2U4EB621ck5HysRV0yu5dybwId/wk3PhjBEVlMOtn6bVeVbHCJcBFgHLX
GxcREHXMtk0uXmEDbS2MdjRk0IYuB7LNHeq8ZGT4v0Ulj6df+lQlFuSYgFaFt3M5YkHsEX2JSuge
uNiwe4TzOsHB48m13PTwS7bsq60vGl4lHxAjcRF+kqci5lgBePZecJKFXY17cp5vTVmz4I93bMPM
ISAafOgLP0dJ5tR6qDD8l3whL4iMNXF92iyYdG5RZIyz6pFppYvvP3r+CvpqsvJETo2tkuJyuPIF
q9gfYAf33t+hkTCVNWkE7cvjHNfuyqDXzrD68Iym+HZWyfxFnwckDOQsawEnY3regIGSySajd//d
zDbYMEi6woR9xAKFFbxxMUvZX8m70xV96e/0bj9qvIrpCJ8fXyNs2UFDoxTKHINtUp9a5D3HfwCz
S+uYOCsdnEDguFH17WyIvb0FcGp4GBnm7HlPoL1TRPjIRVDFvl/asDRNlIAQZmesexfV8vAODr61
c0hQWUlbYzm7D2AYF1PRqlo8axlcSF3IgZzQ2IypVYWhbwkb9DKJwsZMJqjwhCrEdrYngIS8GlkO
1jDb06fV99K6cOuPrpPl+cn+k+a8FwclVn40qvuirTC+N6Ld+oAsdUSV7saM0IYVr+4IW8VrMuGt
vNks1McRTT3E5Bvkz4uDI1sbeZAyJoR1+h7xCRSN3PDjak8uPXjDBouWXA2zocME9vsFawF4H3/o
TOPHZ/bYULoxWz8F0vuzcrQFJrBH8kNV6+YMPaGnYbCxXRMUvPL4WI1be3PdRDndQp45LwJ/y/3i
FbSRLXNPQ0/sR3i+REVhALlWdNgv9ZJ8WckHlU1u8lgxA75pEZnYW/+TF6S3Q3844xk677V08xyX
PSvjBGkNajzo2qo1qNzvgABeRbMV603wS0edJUTaly6yesHFLnTh/C636LSnVGm5OWZAGBDKUiN1
T2AZZE3j3+rDsX1WgExIj/Xu+4jU5MWQ8nI2xa/XaWNGqnnYA5lLXWYxstsOABwAvQv8Z5HVPmAC
T/NPp1Nb2TTKY9oBtFzN3wHBarbKQTrV0Vw3xzMJ0jOfrJXy3UZnZvIc9DFXa6FjFnh5Cvi+yXgo
1gt2SwodxVIEucXVksusuP817rYrkDS73biZO5FW4PCQqzBogonNFk+U17Wqpsm/6LBhpfjeAiua
xBmbhWifyCIZUjGg/p3i1N7hCpChXQcmV/1Dq0dr/EhOT/KcMNe/Ur55HRvT4DGwXwfzo46yZeNE
6NZsrE0/HdPPT493N7+8S2RgrbLSwLQ+wT9FQ6PbiCe+qnq/sRD54BIIbJfBn/OaogRrbgabrPsF
DMVVtiMphHV4HWHjla9e2wWRrC0mnBKN7lztRTM3ZVxI9JGb0ALm74bWKSm7hUfOLCnwriROLZf2
81l0gXO+2TJzVMJVNxbwDdfK4jRiIud/9S56aOTy61tBYPXzOC2Vq+lm3tr8QBQC1KEK5rtgRG4+
BG4fbYOI2/RevF0X2AyOEz86ql+3YV373zLFwmidd0Wn4+9EQdKaL5N5iNtzZ4VwfQjMaNCknGee
Ne5W7pa+Tiy9OTSyrz47s7hIudDjq2/dd7ZRJ5+++BfOBBbkGXNiYnD2Iy1eANKdHpRaiqh/0NE+
7/CgGF0YDpfIu6nCO7/G7gC7CKVQuXzEufrqwS3PEzHYIsimzuVKPaKfGp07Q+WZXDGSRIEV/9m+
auZAeNf6QBbxZOdm3DdxsUXccuNlGvlelruavJZdBoidfjXkY47TQk4lLouEajBecR7NI2H3lVSk
KFa2+5eC3ENYBvLYdrE1pvxgbJW1RyilPw0UcrGBoG3tZSfuNDYWN/EjM7ooC6UlAm0ELqnPpPM3
wWriNH6kMQfBPjQZxSS5R6O/PMVYiWD7SEkgyXm74ZIQNlWhXRbN+9qvwDYyspsNVeyZWucm2FZl
oKo8YvkjTYrkquyx3Up50747n3lRaY7tLwwhvmcf2F0MWWTih4WsETemFE1jeQAaknSgyn0ojONz
Z+eoOTIgkvbexaJxQoq2hwraIxKH55TrNzSsWV5zjVjErhuUnpoqkDk78P9pXhAQPXAEDitBS194
vS4loHt8uEaZwgiYmubswHuE6wUYAR1xiHCukM2rKpmksyc61kJJuNgAnwmcKXq4FQOwFdll2GZB
GF9R7Bq0D/CWdbZeC+0xLGsbfbxG7vwignsIQB3LfJMy2JZzioc6YfNkXzdBN6Zl50m0gQYbC+vw
wtRY6GgsZ2c+e7Lr9hoQMHlkpj73ud+EdEvAYY1AeDOMiLsKKiFGE2XeKg99I4X1IlEPEBeP7LgQ
5FHkEEDuE7JXQiTBhIgSbIdSXPZwNxi9xO4pdeCJ4/WJa8zF17JNgiEELLaN6eqIBaWhVCggPNUd
eBnHLxo5dVKeXRLywHwSAKw9v5EaHU0wQiJe7ME+7HTKsKzvyyYu8qEDTouXzAWkZrZ+2av4A8K2
we+DN5/32KRJvd/lktirthNeH4bIkR4ZmZMeEoy/Z0PG4+M3yY1zkRaViAdZgrBnD5z3278PRQ/B
BjlB62OGB1NlmzybiOwMB03VEfbrGizjEA9VjmEFx1bTg0WFZgslReclw5FUSh6HEQrPn4caI50c
M/fI0zb5syTeMwtqvbSIVeXgtPSUg+TgG4MtUnpFAcqJaAatcuxbK+FlqmsIoTxOhs2PSlkkObaf
i3kovNVVPYbmUtCiSeGsNm/pTozuRGuMMzzyWiQUtwtZDLmcaiPyNxrHqrldpwBD+C5yPXUfhhyb
QNSzFLkwjqlLYc9qPZwjVIJvUl8vbK5y2Z8eDSS0b9NQzZKP8P3nn7QQdVDi8mWaQDsWUrB4wysY
ib0X8k5x8kXMcreWBykhJMICLjrlIPbUMwjeWDv/9VDknAZVQSVMz2iRVKlSep8aM6p+vjUB20Bt
/dHrNxE950F78Fg3qlSCddujxnlOa05NUzmjgnZv29f8G61u8TgULkE5bclVXaMl1qobkxxFqdMt
lzb2GnhKk0HZq/Q9/TQRA1hAoomMMd9EIWeJLeNJ03sntlAVvBZyKi5PTIRYkiX0hENI/dKVZp/N
lwP2VJX8TajdLkWB7fJ+C2ZX0qKdY/Tehj3Gg5CrKV3WR2uSx32ht6Wph9d03uENIlrfR8um09Mn
QMOn8cZf7IKPQDvD6LzgzaC9RbDxZGD5VlNX8KO1fd6VwxP1GGLFdbMq7A2m8lWXnf0WK0T7iWqo
nEwcnyC+owVcq2ZrxXQQCTAEfg13M66HeX0BX7eJWRrORl1wnNsb4/vIf9wmZIqd0COCkDO8DI1f
KnqK24nKvAt+wVoPLcso+5xA6pk07oyh8s+CLSINhCUwm7g3Dscl35u27bJKHPkXBWoU0JOXy5FU
o1eyIy7yyV2HXDSgSUdHkTChHScjOTcdC0vqwuop5KW2y1LitE+F2v6Rpe1h7L4GxV9BBzvHiJtP
Y86VtjbWs5zs3pCj7koB6FgBKZ5zCVIx1kV30WcpiMUWSkgq5/hpOAmbv3lGJ8TQdXa5aYLSKuep
cWp2sIN8ZpwFhnY3ye7mv8QnRYOfJXxOer77EsuSPza7rXvSRnij8IWTn3dACKN/OLVQFQGPwzqW
HY7g0Dz82oyyap9a0wf81dWMbjF01q3OTB90VLJLKfXysC7rYXVhEXaQkgHh3ptv9qz859LkabqQ
o1sAehQLI0/UB81g10WYF5wO3K1+CcLKbEonyg/wCSRCSQY4oIE5AyEdtWv1m5syw3eo+3DmyEEL
ck6deoZsHNfp+4ZUd4eLukdaA6pCnkIHe5GTUBAlxyyEvKN2wUW+0dHy5i2310l3e80Ymqrypwiw
G+IQQHjxUBnDFaXXVAYU3NLgGy4WdAp541plb6xsTOkOmU6LrTAOoGp0ZRyLANHcPWSkBfl/aYo4
cHO1H9odAsf7IvU3UJl6asMRT/EzZHkfurfkY/xVaWq8K7CHxR2tTWp2kyejJ+mzCUAW6xBMGE2n
vHdY6xMz2Bu6okzmmq9jH6tgfg2ZKQP+qP6cRB7iye28XQCHjy0NnmGTUZ0PZhzZjjjtzzRvnXo/
t57WIwbcPkJ21FqRBKn3PoLzphXenUB7reFkvvlqwkgPAi0NAZ+wMMSxCTBuauDy2oUMwsBV5XMk
z/vzBZvQp1I62UbaEKHG/FGb3v/69Zl3WyKd3az9aQb9amXt1F1Q1bcXMayzpGWwkq/TA+EgiO7+
cZ1Bk7F8mIivYg9CxoGPkw+KaEfRs6DzgQmOBn6XWib1Qz5QELW/CIs9+vtd+VkzT+e2pBXrP1wx
AzKMgZWxyjuaxVghRKy7zWi7FkVc/6YiNCON7Swa4ZEUyJPB+c+EyBHtzrcl5cq3yv6+OCSpWU/p
ZSlYXADSpUKJwhZ96M9GkaY8wVkNUSAuGuXE/ZXby42uNze8lmoWO1w67ZrtFae92PPhTgu6uLD9
5sGv6DqfssKbrA8U9pwSyoaxdJQy+WZMQwP6AXMO2M+8+eOXG4T0xl+WE3mOeH/2Zs4s4M7V+5cu
r83yiaV+pHvHXa0OEBt9Po4rpIwa/haxccdFc3+W6cH91PjX+MAOUlX8khxuB84vAU+7vIPfVIcL
tgkLARa0HSkLYU1r1Wf/mB/nqKjIWopVB8IdRRrcGddzz88AihIHdB0q6Uei4tG9Ti5GxidqafXm
HC32inoIK29+t4EurcbUvZkiltMBNlD+rlCN6nYDVJQrE4DgW3GdRDj0zyEuW+kR7M9NIcWZQypy
s6fdNpP7xHRVLV/mUVPsyIrbat3MzKIXHeIgMFfbfGz66cUdwbRlmAiFGsZ0N1A5XOKyh70pNQVj
zfJ5HcNrNGBfOZLTjRpxDzyhxuO2tjQSx5GRQBoYjpGPhcp7PDkYamviz3eMla9A6XWKIOw77VNE
wZr1tqGCAy69ZKA0CT5GKDYrZLC+47hYcSKb0FNQFZlysLhX7BX370NGoB+5Cne0b6JZwzTprK+Z
befRHiyrls28BJtqY4LRFz+3+ZOO37oqVlSX8NodagatL5/fwv/tuTPneNyEGZKjEYJiI1Cafh9x
7/GsStu2jat0ZG7OEAQGaEOI0jXrJizXXZw08oD2Da02IfCIIeQdUJo4Qysf7WoFRpebdkmRvmIJ
1NG/fUDbmOP8ebrzthk26Fxgo+jHXTlPzW4E6b/H3ZMZ4/X0hIy5+nxv/S0062iEEtZpmMKocALv
oVlF25J+MZzGPUPPDs8bsIn7yifddYFkVTDIEt4GrAY7YeZFhrxJJRzaeS7lHkVVPezMDG6qrQca
SK7Cz/O+9i040qeaGokArfkjpGaeJ1/MinyjSfTqVACICX0gAqYiFMQfxJVB6LNRMNR3lY0ZZarS
Kx1b9xayXXw/Crx9Kkw3+bXGV7SAFN2g+jDxJqRZE6lNDkOY6iWml7sZjx4B6Y50NMyWxdZ1Y/dr
2PyI95VzFsrqK099dBZDQXk8ietNbctPIJZhOf+EMDqOnLrqy/KyKUnojcC3DX0fWdpduJsGsDIU
O3SzeFED57zolpTVtyKvHbHWjON+oPwarG+6Z3VUtF5XX7H0we89eQVpJTQLPJSCtodZvtfYrwBr
I8kPrWa2k4LtjproxKt7Tst9XMe3GBuKNVtEMEW0Zm5SreoL6pgTBZCAtbSQGZd52g45F9DrkNju
nxZ9XLF+gryn9hnYnnJd53fdg/fJ0yfK6LD7PXES5v7FIO4fPYwduLDYhf6vRFRIiPFWngtYKfko
5jT+yDOjc2r6d1zlmVpzzvhjLbwgZeGBi0pAhZFzipvDKR554CXmq/tPCiLIS6V1enDEvd2JQNu/
9dvyCKMxz85eDV+AS2iGH0M3sODRBAEH+SKrX6GR0jXfByTll5/D07Am92OYM7ezV103isv2iYPS
gOMdckBQKb3NzjXEF8vUGLz6aUcHmvNFdsDxF/TXnpI3GrnAhtLsRvBTWgq70y1bsk0PSNkAxGUq
wEJt2UMlJp+lOAJvIkoNFtUoE3uC9xWcEgE1bWSuJhjXUF7eWQUzm/T80UT8X8zJ1x6b6H67XbN/
eCYHHWZ3k55iqwKNUTP1t5TBqm31TKwEniu6FgNPRQWJoHhW4v6BNt+XPax5noxaRpPjFCENrKq5
aaUmQiBpNSEgWg6XHMET9mVEJU9zlwLG0k9P2OlraAPcrRMkz3y7kRgxjyXqleEf9dfHvZNkhMt1
LNRC9YkeDenw4xw10jy69DFjeqq3IWVERho6FaMWGiPdSnBuqBQmGEO2Ut5aUq4i37P0VAnNxmrN
9TWLTLnz5o0sf/kFssegqaP8xYAHuBYsutQ7GAErR7a/mNgwmYhiiAfMU6+xrG/u5uz6GTMeVwlL
GebnQLKYh4wmO8AkBTNT/mSt7V7oGPl8nZBI1VBvbUDHAHONit0tkU6tPfqaShKHQ9SZ9VgPh8Ia
PkMEmpH9/jEL8K1iDB5w60LhawGzo/kT36XWOqb63+uO8KMYUvuoNQikeEfKH4mwKsSgCjCwlxES
kh2aEmXs9Qazvas2whzfRjbXr2f5Gjs1XaB7UJDR3tp4VrdAeiWLEXoTeO7H0uZptpoBQ5q89vBv
3Va5uczLOP2z5iZrk5CZTG+gg3rayemHDJiEw/U8RhRCtoR5jh6S0k3TL5ClASI5T/H8F9i51QRp
hEcesaRoAfmwg/onf9+GKKrWvqQTnZvEmEerVglzvnDWORB6BJ9/+BqwHdYYa54XXChgPHTYEIoP
RyTBdXaNYNn2liWMuS1cvoZrXDtLNciRCyJevGOFl7L23oZ7unSk9YAy6/TiFmsklDBegV+NfcM4
VMpxXF/JYlqSBv6udEnC3vgEjeg/ym0IUBtk18EiKjdesMup9obrjMG7Mvswp/WlkAKlgskEwgfI
kJKFsOt94OL4l7Fb1M2Rrth/aj66lwlzzC3RiHPryG0Kc5idBqGBIXR5PlZq77MY6Nb6vcN3EslO
SRa7DLgv2uJ/MIPiECN5J7WSp5z+HaJurv0FvTQz+P3NHevslS7fh/5ZoJdJ3jwWMuXIylY1ztC/
IZBeDtXYfFJZPr68Cl1EQEwidXCYD82M5zBYrwHaWr7H5Ru9bJm7nnaKYyrT2S4XaL99Bl+gbqzh
eErnarPSeMUAOHArJ9JDdZ6QoCWNYRX8q3mfkaWUOAXe/IULU1smiHJQGxxbtMK+2CPEQjBUpHeI
2IHiPM4sTIVJqALY9MXlHQt9sTidPY2+Bb08wrJzRqp/j2d/KwmHWb/GXd67rr27qgDN7hYPh+dv
vt/qcPrmsmai2fJDBWd9VEp026TkVr5aPyeiGDbjwSemoQkYglFA1XxUlq1azo4njFzVTrsYmgBF
VCZv4IrqYh1/Hh7kjqmE2Se2k9siPcMkqQMcQbpOGSbTqRn/no4MFjWNjSqtULVAmvlIUMGE54mR
7enn3j/faBx6Incm97/yWM4Lpj9R+TuySClTyzAPFq0NRjfAtlXf+1YBR6rTuf9SaLDxGx2EZroV
dFHKLoNvNMNuQCVePJ6y3JDJnzRAYecBzAyfLH6n4QTcvTej0WSAr04GoRKv/S3K/PRWTeL7Eon5
pBdsefIUIrw1VCFU38zr/wYjFk0JweNgU+Jo1hpHgqZO1A62ifc66VNnGzaxasVsAgLhmuq2CAyX
2GiXc8Smkvhyf2LGyX0L6W7jaKsbFDGY+pzKmeRhx5wa0+Kp7xsMRNhQM5ng+ETniZ0YqisIutAO
iInEyIOdbSTh4Q0/wFPzEXbnhMGhnfp2VazeODc5G+IKh5EVPqZN2oZCVm3Sj++S9C+VYVnoCHz2
mONAFR/xtnrh0fX3O80tgrB/flIljyTMWuIm74pySxjpWwKKd48jorN/XGIZOMv3kfeAp+ThO3bh
UH01QH3WK+Os+kLGElTpNGGn3NI4KVbdGWhj0fa1G76OP+7BT0dU4Crbxn70uUI2ee4y+NHJOYo8
BCC3lAnfJxeuZgUMtC0l2iH+jTheg9/PFU9bxat7yF1HbD4ysmupnSNbBqczKLnxrcqOKK6tPlfB
UqPJ9JCIhDngRkIP3CvGeBC6mFGNC7dsK3d14trlQ6TgdTWdsWxtnIrzffAKoFJyHX1FwxD1Y9Fc
zQtTvEC6bpvw8lcTWpX+GKxqG1gUEtxV5vxwHmLH5topNv18QppBX7PWSVvPy6PiJOLcn9vx2TnO
xTr274hgSViZELw7E9tR4m81bg4tERJ+rzVkTiRidR1aKmpgZbp7JbNb2proE+FBahrGjJrmB7PF
O0k+7CDm/6/sVNCwvkYXK/CmKAm49imhpWuv3DrBJZnULHVcqWLiugxc3lLc2y6fD21A97/pUu00
3cUnRGTs6CzJn0iV3v1x5GJpv1vsUUylUKt3DNwMmy3Q7Ga4ADL5qUCnIlxD0hO2srPvFZNT0qbF
4caRZ7K/PpWQCaJQXts4ievbNlUX+tjJ4ZNh5tqZd/hNT7i58OkU7hT6rjyPQUNbcwfw0vSbhvgh
H8EVt53U8qia+uvyNF6UN0NfXvI8UAxrgRT1CxidycxPTwykmXAUT8R0LUTop6FmAKv5f8xir9uk
deYEFsda/CUHBhmxEGUhF+KtiyvYMwMvRq8TppgPE4TV+FIuOZaGa7NvQGpd2+OwPoRTDezgc3ty
LmqXUFBMFNaMtKIw1yVLpVVjNXamfczDdkOF16GZc8iTOzSy5A4zGBHa7DrkHTsjJZwMxuNtyVj0
5F8wXeUmQ5ocZqxO3iMvniyHa17cUsfCIjvzuq2NH+Cj0DCb+AZa3drfAd30+MQ1wYA/aG/nvonn
N5DkDLTkeI/wve7nL+tWadgaatZzx3TwA3vbyfPKQx+SZaTlHtmqGXGVdII8InyLGRUuzQl7bMrG
8i99bYjrklb5KszBNO+t6WKGQAPKMZv5TxsGFdaLOB+wf3myVPYt70SKCwf8hO9OWhWbz8q4ycWE
mF7ZIGfW4hJSHa6mh6gPHuI3zQT4ER55nramShuz9Nlds0HL9Wy5uwRCVGJ9LdQ305WCZAw34e/U
uupbT7lxB3In/DvQqsu15r1vbTLAhIXc1q/2ywTH4TalHb9isXw5TPuemOYPi8fGWKPQ+xjt8HK0
RszAl8CJXqMDaQccIPns+EyzZKjS1y00Bv9a+ngv17sQlCCybUht7KMdIPqulKIIkPncw3MB2gXJ
3G6ET6qhxd5132JVmG2oPV9VW3tqrWG6wLnFCFVNT3c3ysI9Tvlla0TFHp9zT+QdjEu6wCgfYFEB
mccNT7MpIAC/KBHOwNBvwRzPgCamFCMkI0xJ7ipL6f5zeJ1nAwHuYLiHUrPD6RdRzeOGPebO9C71
2KciWjJKdmNdqMqmY2GMjtWjUzUlip5/1OWCTfsuW7KtkBmJgZuARu3NvmqEqtbKrVV7VabNXmWr
7nZCzw0BLMMRRKIMO6+R8q47KvYmmdE64GdHcUEI3mvoqSwEo59g0dDvKEk75w0T7y7zmZeqjn0w
JOnrKkJoLfBwGz9lBf6RgHltt6Im7MbHWcNYZ/y5keWbBbblrGJJmXBE+VthPBFwhJpfWntXLuSC
Z/qp9RugwZj3pfcyQSYY6nT8OS82Mw/6Pl5pnkAco2DPuQH/MHzCbL/lC9yZT4KMuftWjKm9hCui
4qXImTBt3+8EVpOe//OuGtgFeGuUGTAhFsLbtRILLK6GtJOUa4MN+1rIbZl3F2SOsRM63qewydS+
jr4H+DrqhXdm3Ic76s8s3uxmGs4RKbwuONIxptZkQRqmAL+lrxQueSnjxbb1p7ZH6B3TAMp9Tl/+
u/Zin8/5uuv8PVCxn5+VzQPaWHNEvP46lwZpq6WQKh13raovP75t8kLTFUJ+vhBzCrHmodL658+u
oa94T6bIsd+cYPaT1apphDIT3PJarXB54dryxUk11EltYWr/dUjqpjc9/bJ0SP11rdVMHII3BvjY
Us83emQ6LoZGttOTDKPgFVhB4CGlQb7yF99KWziU8w6KNIT0pH051sBLH4cvdZY6ndth8M8HcYLK
Fgjmpk3GrYpGCn2tlWuf79fYjtdy9U0IsqzzgK6nsIsnvMCw8fl78Wt6FeAwFCbGdFhPWyu2c/6R
SjKWa4MMgVMbqeP7Fv6r9Bx4PY6JrlRE3L9PNaKNOATM70q1zfTa/LjgsvSBmJD2HYTLwsARXeXM
A4tK/4w9wJKNzbs09ifY2pISOLnS379PRNo6TMiBRtpsXnhpP/3dZ5JUsgb7ayIWM3gK9Q36EyG2
iaP5lOdsm3Qa3Kp28bqwGXWmLq61XT/krivYxO+mkPp/DjUvh5lHwCRQGtrQZqdopA1f9tZUhHg4
j2WQAufnwUTu0FtipZLoDos3qkS7VlBy3SBzpTvPSWO+ekrAjo6SzOh3oEk52ovMMbD9Cqct1Td0
srK5VrDpmdg54iuNUlOmMoibRQnHXYY7G1o6FuavlAkDsgiJhTeNhtUxB6ZjSJ52Xyh2qaEU0e2s
9qKF+IPiSWpkXTAF59x/b1vAZ04BY1bY1/N242fOytHGFw8zUwJDwjn28W0qXtbChEztHn/x+O0C
WSmOAYzJ0n1qzQY9YyRaEybRviH8x2kNuTAbelZpWnjk1Q0/dDFeC4ldRQgfU5LJgUpHFDOoBRwD
2lbNHAQik3rOWR7gl1S/yqTJGl1zwimaI9cSMiuGIKhZHNtM8P6idaMnScOBprTZ4nXeDUcQX7tv
wnCA1gOXT6DT52bb0cU5Qriuqu3wo5VkO6jaqwF1n6CJ8u9jiis7u0Ji2L5YUb4a2kWajCAfsgQM
y3nC6COxs9zcXT1GPmwSXmLs+ZdlfBw02vqYzejKX+mFQbzWS1EsolaeQx34cqKJMTtoUP/oY79P
3IborQwDn/4dFYzIGxQtkkN5qvKlKfhDnLzJ96WB3a3t8XOGTbHATls3n6cqNAeaERCPRI+M9Br4
Xfj7Mj+Trr1utjRxQFNcjk0+Fp9DbtMbNLXrI5LxJLN5JBdknLqJ4TRc1BJhUCWfTtqjzRlOvLUf
3DJl0/nnIkL0x+ZBJVzBt/dz5RCoeTAqDXM0gI/oqd5Pa5+VAr64kw699gUIAxr7rwnD8x+qynT0
aHt0Uso4smEOQr0QR3yfq3nTANtjMkMOIgODswXrAETFKmiobhSrnt6b26MyGIOc2PUtsTtB6mUr
ipJPBIXC7+1U31cAIxXMXYp8tKKD9PTRxaUJXc4dgRWrcDWZdjFW/1+jKUAsEmlyqdwOmsQneEwt
z5hooE/qa+7XYcJg82Vd1dWKyrnmPraH1ZrRI81k2ouFHJoESNCWRXunH6cTBhnNs0dx6M/GL0vA
5Y9aC8vJHx6IUGai76gda8SCyWtLJ51BbqYnAhcmQSJBsV9hKdMElISkeZ9jTQGCvWBudJfqn2UH
7qj1vcQQ5l6FwS3n4d0uH+qmKFPAxKHbDb8AtmM+upymqyRfTGWe5XlK4ZGGUUOzwo6B+VAdtwZF
KSPWEHcTby63SS66UqBZE02Kpw2v+KVL92TFsfLi2xZtHQpRzZbPpwQ7la9Axky1xV++WwtkPlVm
0JxzFy6570mkHf6GbfGz3ceUj48jzaj0cl2Fhv8Lm+UuxR9Z6YRkdWVWPmzyCrhSvR5Y+gvWRg7i
dgpTfDoHxdrB91Soq86GUkwrMo3wHlLoqLbLsn2f6TY3yg40AY5Akt4lE5wBR+LCnEn/VuLVVzwh
N6IXYmkaVmeofmBY5Dd0sfgcaBxeTT2PeT9PvQN3c39dtCXYL8IZ9GvsXh5odokaiTD01sU6nHXL
lCsJL777R1cIKBH1QeV3p2WK/A6yn0IsbWOngRa0jZ3evmjQrWML4x2aCPYP62kW0wQmMM8aEqyg
65OAL1pQXwxx/cckvnDYOWJrNykZhIeMcUCVHBot2Fgtg1/hyOhmM9kKYqMxCz/l94gqDyBgQY6h
3f/0L1KogOA1uPYwmtW7k1OhswIlUwzKTYvAGA51J0M6RDIFbF3PQoR4E40PHqbu+f9Ai/Gxw+Qx
bxkuso2p9R/57uSxBf7VflH6uvs/eDYLmU42nelhlUqh0R6UCh9hpypTfGgC0G5yOpoG+FqdqFHp
qNlAd4Ubj9knrgGFf1dxd+qntMw5iTbBnPkotxcLtRxzusAuQSs1/Fvxr1auSRfaqRxJrOfZjClx
6Hxx28BDg/xG9FL8zv5ky5imQ8ocgbhqLxoH0hdPZr3xVNWVPUll2Og3OElEzuxgMpDsiVrilAo8
Y1KXaaoBQu/WgIBXFsxicodPLikrkWd1yD5KcM2MbcYx9ib2U4Yvm8S573fgLj73nmCnqQhU2YIT
gVzr2GUEE3aXnE/u5TTVz15SIk+B5bKrw/t4kM2oxQnNIwdoJBnwXvO5D7VKTQD0TgriWnZte/kp
dKzEJuTcto4Ni/6Ni2LJedFQgj6LrgQWe3tM6NK4srF1F2uh/NmUS+TsuOxKL/HDiePGNDwZPIV4
u2zPLmcVffxvMgCpWZzJKJUuFVv82VlzVqWSmo0BmH4pId85X018CtmbPWWQHbU+FZGR3DF19xIi
N+jtQ00CGXOSK3UBAPo7Cp1pdAtGjlzXLNJhD37PTa/Ecv1ca5EOLMWEhQFXjHfjbPR7RaRp+AXX
KDfmuFSlVQukTjF1gUFCU2t5otOCI+aMHRawXof9Vu7Ly4sUQ/21X8fRdJHbAQgjhkKa5tQfMbN8
7dmwp1eQsmJVKJAxmecNEX8iNRL5k27lSOtDQYZ/sKjdxc4D6HNPtGqtdwSwoinCn1f/AHtNK6SZ
eJ4GrPjSTVrb4H9gEoil68jqFhJG9lX2uDCg+gFwjiaGJkKSRR5D68HDirLdogec9B9RHLNDrddp
RkOLH+VrOJy5OKA2H3hdZJPt9MXtbp4K/wD2RYLN+zFrGmNgjRGWeAosXgaDTM3NWzxcQmQv37BC
dIInYidoSoPlUREWmo65qcx1y+KyDwzlP6n692MJpb1a/BaYBHOTwOdQLg/cD9fuFL8uY0FV9JpT
gtQsZZK0/O4Rajkkvp2xawAo+v3mMbvvJgHrR1IVRJbJM1DaYAe0do2yjUVhC1/vx1E028fVYqV3
zB8G1kBgv5T4NNm2uaC0aXaBk1wyxgZYL2UKfoqdnINMxvamui6ZicqCWVFq6qz7Q+nJQ5igR4Fs
dAaLjRN8M67HHiJBK9jWZ/e0T8+e8NNLMNO2nGGCAJpZa+BxwPyEuAc81/2N1Y32LW9VrwW2L6aD
31Po8VZUk2f9YdJ5YYQ5ZjeZ1UcYv0i/tScfGiANYKx66XscimGcTVh7Mo2Nlt/aBsFR2ufqGZyh
yZZwjfwQO0HVpyH4YMFgm1Lm720AHsDR2d16xOU25vVKA08Mz35S61GswtIMY8hgVfsomHasJb5Q
Bw+jcjxTdc2nkxinsRRIJ/BNTYvuLdWH7mUMy83rV3jNYNp4cP5Pat9pWwEwZ9wkOOF6mx2+M4y9
vbTFGmkExoHWzlFQBJUJg3OCiTRyK32s3JyyAU8vLEBi/+mSVtB5tC6+fxVQAhqM5U4K8QuWrnK7
Eff6P9G0hQn9DhQk94NvEzJsuv5PULg3cnXhMRY192+5TdTT7cEwGxqRTLe4ztttYMqkLwwo8XAt
atMGeLkpTD5d5nadnEdwDN0+9Ck7PaYABWazSmvxJTAcFj8e8JNybs+G2UJBLoQGS+KWI0Rz7AvJ
6+kPgIcu8XkFgaiDJ+Twr/5GrWmYqJCWKu3DvKrcuDt47JjHSZsdPGtpkR/d2iW168e5BOFqP4iB
pT3HRqeM+tl2lp1PSm87oFsVquMPd76QA5bFhi/3iCY6qNpKT39FDL2lSFRuIsvYkqLtkEym66he
3HR61O1rcbrH/g/RnDpWEC1srkUWyN0RtT+Vp2D7lI60DUH44rG5kUOOFWyC3iJ8AY+MTvrAftOI
q24NlIKabhdpMakah0PyXtdK5FhoRGD48c1cUXC5Vm6XFtPqfVT6sDbinyn9OAy+022RlLsaLJJl
oiTkGVGDxevgqf1vuKArAhZ0SxUyzTN59iWD/TVP0wQR+dQay9yGkC8T6nn9a3A/DS1quIDIikUJ
cmgBm1VZ3beEt/j0pDdlEIiqTfsEBgZ4xFy1bmhgV974AbzOiMWs+xywv1cRUrXdOXesYLXAhA4+
qLHLQy4+88KMDqU0SGTwOKiCVbz/hbc2n7NhlOUxrmIwlFLd5xPgZzNX4fnI3bTvHr1qZYRzN8qz
y50V8u+2vvIf6SZiNgCRJwm3ON2a4Yvv0u/CkQAkIi/GKWf/JkXwHyfUFeFVp60Ff4uAX1uHdwNM
Dy9Q+AHbZgm5s0qN+qs8keiOje5Gm8LgH7sod1j2Tiep5pm0gdNR0LwNQ0afkrYVaT50l92qiln+
O3noW0lwZ9FMB3NMeF2zfiC0zGOBKDchdEEX5+/rUqOjgntwJ3TArCsvkQiJ+1XV79tW8pksjovR
URs5xTlxXsr6yItjIjW+ncnaz/B5CqODs9J7vzJG888v2EvivnXr1U4U2atqRqP+KW+sCVdaz45h
y5tMGu8Cz8veWQgJTL1NX7t0lNoBOw2gW3SJCCe3UcsyrpYcOLIGh7pHTlgEcerywdHwO+u8uuPG
z2GZGGprsxfD2uT+zUYf28D+StFrq96pPwnnJej1NN/oBveEj6jqL8bdwVFvygUQO2caNmMTKUWE
RbVjQGYMzsnjJJTyDU+JGyluwsaljl63SUtheMiDR8LKgmLPKDEC+XXAC2w2g3bIvMIi/J3dugcg
lWyBuBwxuxcISViUJ8oRNbp10Fpi1937AWP55nPBHqpHj5kmP06iUq/DZ9mQLHj2igCAU6K3tSnO
kVExBLXBQPGsY/6ZlrllUFDj5kjSKcaCTv8wg6qCQHs48cXn/febz1sVwXvhf6l3TqGLrq8jGZv0
oJqyvc6jqHO8SWNEfXvukQKJ7zDAqrW4J6EomA1Z9xZqXGczGJ7maa30uMrA13IjTjZOrMMc09va
GOP/CB+4/4duGStcugZa6KqdjSo+UD2q7le6EoJ0VdomEi3bE0yjwKBxhT9ukX7TuCB4co03XBrZ
SObWpuOdYtmgMtUBUj0BwILPNRzvxRuxBen/xyoU5O6ANKUe0Z6ZtWzFxzVKxG0XrWe9+HObtSvt
sVt9updkqNPDY6KWQKPU8YCwl78dbmGZ3+cDiAVrQfVtGmZZ6f6/JfL6QZvEKRJ9E5m0v1KO6e5N
O8jEfUk0/NtVh9BK+VNhbe8svUpG6Ju3CcVn2R/LxGbtbrmLXI1ah998YevODfULXf/naKOxLsp4
Qms3TD94j8BLzVspHwSO6IGYkRmoKw2MAQ2cmuY5oOUOpZcOBoamSoPMsqtaOiwb8/3y8m9OYNxY
+Bhqd7VImyKvbFX21utoMYrb63MsS7DDSXvEy14IrWYUrnistzjdbUWKxzHJd8TKwAwX+6Ufluxa
aJeN21fkU/85Da9DcegropnP8xEI7GT9ldPMgFS24DN7MGcxFuzAnLSFIwTpo0fVZg5QJ2im1n/P
zktyzbGFH+z/i6Wqiwqr8cI3RmdVXaaQzbdJ3X089FkdB7tsTOXDhJux5A/ktMtb8LKDWxpw/OHs
Ts6Q5Fwsvvw/BmVAXZfSVx1xt5V54FXMzXOQjo5WUZjr+VoI/QOpZnd2q55chGWUCUkVscKsNaWv
juRGUEbCAbIBwgUkVfkVqVoT9npsS+YXMQxPsyOyh2mYVmBdxT5GcFWcKdsUrsTeq63+2fBogorQ
pEjume8IqzdHVjU3U6yCLT/usdUtvA2l2frhRL+SPi3khH9m9Fl3M8oIOgzslRu/ZcybKhE/Bprh
+5GQCDkhlwzh2jxLmYGcHtSpuncksjFit766It3aoejlAT0NdwBdLVNg5bMVBZJ7mj4nFQjZyXtJ
4hCVibJfU94ZjpaXCowc8BY+m15IH5j2oRiuBk4XXLcwU4nZPFLbWPBcsdqHilfGAssGz7lD9U3S
SUMxc1kZgxCQMylpevVjyXAnBUMhWdBSvGLP9InKZ2J79VggbLfTYomNf3L0fiB2cmxZwKREEK4y
RxkMYo20QDDYuWm61j0GEFVb1JLc7fZxNH9Dp8fnzKi3WJgM+tdrPRnXS+T0iop++QfuJy/P8zCb
dA/wh+MC+aOjJNnDxiW/8wgfOZg1e9usA1+/8sGIYNZnCp10QoGKp/7YuUSOQqfm0BaRjx2WJaq0
i8raSOJkKGH2E2ERjr9aG/dYsAIAqYqzgcQbjIzJ8WobSDDVXYsPi6+zE0xSdzg9MbykHS8IaWsv
2xhMKqqCJBrvLki/h9FPjZh0wpyD2Z8wxgyMDXJzmd76qCK2trnsnm0G15C5c1X0FsLmI5Tgh10l
RXi5KGebPUKvgmPiiVI2hVdwMYzBlPZbQxKxxaXw8oyjz7FF3YYngNgACIiJzC1sdivKrZHPltPn
a8v7OVByPot09AJjLL1lvjyn6IENzsX2FzZ69KWZ6a096NDiHQaZ6yNJsTuoQm+gkw7WzS+TAhM8
PtxncMiB1VKVvswwa/B93zPwn7aHP0I+n3lOCOy5lqJkXcYNLePDyqjaKKOIXFWxVDxzxrqLEKZC
LOYcHMeaPuZwPwui22Kpraq3urBCUOxlC22IAWD7LCxZjyvwzUaoYvAnDttVlx6S2yMBZTix+dRR
0Sv6RTM0s2Y/ju2BCFshpUi1l3WhjTIsqARqysNipoULcGlZtJdjdOkFUVfBopT+Y57FipxloxaK
HtBBeZ0l1mGXgIh/IDYVOLpNf52kGV8SjgTKRM1CU3yxJ5t9RK/ixGsnqVizirqGx7e1XO47Gs26
nF8COW2k2FMmA7+GnmBGNguwXK/ETZRCPwBttN7j/X2R586nzBjV0191L/VVGu+wiHJlATElZaNK
hyJjkYVJgi7ir3kLAwMmRee6jcROsVy9A7d9uyt7p6jpYwwMVC4sIWZiSBJrH42UbTpOZtuO8ELk
Eu+pBzRKQWqmYZ3ajuE+nJ0qsIBTFDuX0Rxrbif1UIOMmOiny3M/YNbpNXg0gqajqlhZY4KmKRfL
TgX+XyNrJa1KrdVg8HMhoYxmBV1VO+b+4m7ke4FzBe7TeoqcyIgKo8D/T9LwyzeCDWGVkyRij7fn
wdeBsPxpRFNplVI5Mqnc7GByZiCiUDo0T8Iuz87liji8yi5wAMUyNqEH6vDMDfay9XP96GsP/o6j
j2F4tBBsYKY7ykKjO1a8gPZeF4UQs+PN5u9E0ssZD6XJG1hcmOIgwXpr1zYSCEOGHUFvpCy0Yg8u
7oZmvllR8Cvy0D3p/aLjNTxE+HvPX5XAZ3I/5McKlm+mqPn/P82z1meigZ7HGS2W2usfLO8WqPHj
BXWSGKAbD5dh0KTcK62M34uoKXqHoqaknloXMEK6yP+I/si9VafNA0wckCnj63alvfvSEnDnJYj1
bb9YYc30c7pAS7mrAAM1+DvbSf0d4F+S5K/i+DZOIRomaOALQ3eLXT2i1PV8WbluJCj6F7T0y7o5
JuH/mOWcqdKDp+dogKCcKNLcBzY1cPjVTqZKVyEsNAcmetZ7Qv/khtV6vmkbfGC3873/xFF77Zcu
F2huTI05SMpLp+yMbCCwkjkZhx+zVADE6WvtcQC+pY8sPAD/D6PiKDioXN3l8Rjq9OuEoegUlc23
kSLhxxxxy/bhCMV2Qxa1EnvHfbfJql/iCCMb+hHQzC5bLtDYmuLV4EhYcBjcqK0yg7ZZ5+VEgXAb
0OtnAtD/sgFuT+TAVUGl2uBIpZ+cCoYAIQ3dc7oIhQDysSVO+WlU2OD+Cy8g3S6uHgnwDCgSSMoa
ElVXFeW+yhsl5ZAP7L5j/+wNaJ3902rLVf1ALIWyXhfpgkio8ExmvXtiPr1m0GkgkdWqOh3wKtJm
xBDVd4FpZrnkDwwAeAuBdMCKkNMlAeDrjvO5Ag2mvPu+FGdBvhmarLQPds14+3byFKBs25vJBxHu
Zc6SyIcPVxPuGx0rKZBQAnIBiGWchRQh/uR+eeNgOeUUKi+N12uMGa07oc29TyOCGlMaQrsebrYX
cHbnJwmYjQ4HbWd45qWtqr25P9mX15RGbgOc8DJgvp+kgtvZmKQeW7NEk+xOaI/OWaiH0oX9VCe1
dXoq9hDp+8ygd39YB+vcaRBeo9X/lFmx5W3K1WQbDrZpScpadDe/pB38WFRLv5JuknKKOXQ771LO
FXqQBvSFrAz/Q4gOkslFAQXiYIHYnZfRAiGwhSS7/AF38FblTr+DMa1oMn1PKw9F2UY5fuOHoWvw
eSLvgjeic9vo5yxHsuZJSD8YGhhvIa8ERIo2+rUN3XvNLWuIip2vrbeoBO76oGD/b3lwQ6CUXMc4
FRVegAN9/sawaEJW+eYoaZMswfozL5d+qmt5ecgxu2hvy4DjOy4883LKewnnIly/8k7rC3h5FAog
7AhKkQOsFKGnJm2HiAZY99sa06nyeuOLv2UFzFDpzgkQcIH2rDsbF+GCjThEAEurkBznHOolVW5m
ZQpQKwlf84CIbuG44Tsx9Uv27vkNAFoyKr5k32H6B8oM9HSeCufmdKlaZTR8a2LesqSdA7tKmZSM
B6WtdkbKErBkvHpNXiEBpNkc5FJUySXOZ5k2am1MdMmQjyC7DOWmuk64aXTGwjZ/m2f02wgMx6S7
zZEBLWVUy5Yc83vj4l3+BVtkycb6rhKMxt+yEq6+ISv3NEj4hyEvvvHGe4c78QpYk1hSfLx7QjKq
AHeISCsIszL+t/rcqiK7cVoSzFXKp4S6RQl/SE2ax2ok9m91TbbEEnsRR9Dv1PoLF/hczZrB05Fa
Xsm1aDXrrSBIEBcQKHUoEYeAXePDPExZjSp1VoVjJKOOR1Sn8JQrjIxaCR92F2X6PKG1yvX1c4ix
iWPo2L4JYMXCoPx7gLVDp9iB5TvFveck0JNuPYoiObBbCRZFRsjLgNAhYwwKW3rbZZHo59w/StPp
DbNyZjEjrUaZ4vNlEkrpspGnutldienV2/5zuycs0i/0LH3nG5IFuaJUCPmPkfT+ZZP9GOUDm43c
gaK8DCGiZb2RMjUSyPAqZDVBVB2refViYfw8TKIGslyku9mP51tPaJfz18cYjCrpdJPxOD0XzEdu
EBYlxQt0avIvvWO7XMYDrAidllXF8k806fn9J+8h99DcRaORSvlIhDnHq8EviijhuDwGPVLfb/s6
J6LBnYtd7b52EEXVr35+PQeYPyp2oPvKSFJch2Tcs4SgPyGryrnwfEpX4tEBkyljVrQ5cgvkZDLn
ZxJWi4Os07776tN8/KSqpOWW95DF8YZHsKoHVbnvrEUsxG6ILHAtsbilDYkVLhxBRosskCHqLGbR
dXyCRRU5BXOjOccLiNeJUxoJ5OlqMLgGpaAGnprXam8IWGy9Y8GjoVTvUggoXjpPvUkWDxXJgreo
APy2RTsH2AUB8AABOazoUmsQ1ZM1c9mPCGNnhW6dkFX6AfJ6oIKN6sqV0zoKRYEGMhQxRiXogpOC
pOU9+y9k6FCeRZbeZeyzmqFW6RtCGh/6OaS+r1Mp20uBcSx+N05iYI2p8wA2Wda53qYYx1a85cb7
zrAnJflMBvNGQf/MO7RoTebZu0lgbtB6dR00cs5UFT1/tfbkdVYeNjYE/KIye+BskQqNzHGonz21
oQr6URULLGsuC5teSGx6+BLubMTplUJkGCLh1T/h6pXlb37O9d3rqyNm/VCkIC05+evXg2qB0rxF
MUavHCK7+2NGst+no/Bvjn6uUD/eM0PW1cFcWfTnVcxu4qxw6y1UBwnwYBw4JJRAWYD5zA9IxTXf
b6oUTWrBoqYWBnnk579pg968skW+efkIVLZAIuKwJRO5EYq+dE9/Yo/tRxbksXpI7838e0YKSgSb
dYaSbG1lgo2riooSDoROuMNioe3PuglgzvCS+QXMbtrLuLUKo0hOkimTuCj5LBpn+BuXjt8oeJ9V
6596Q2lQQ24p7dElWWEnPw1xr6z4gTYjnd43Wmd+q+14d3SKiT+bYEV1eTCyEWh7gTV8vKCzkwp+
WRAF62eJWT52U1D468UNFYHbp1IEomYeifs6ZmDJlShhrNYXo0jfPqUM5ZG4js+U7/zktsWPFo1g
Ct9u6d491ZXU5Kq7kmdNM/bE3HiAf3UNKfLbxYKVCItwk0x1fCDQt+18C1/wXc5gVupTeqX8GyOY
g5J0c/X5BjEk6dBVTWW3oJzNqzcgnJvMLmBOKdbE+HHguG1kNqqTc5EjxEwck5bWgKo8o/Y+x/Zw
VkvhiF8Yo0yRDbMdAsMUaSH3nN1v2UGtVm5a2gs/ERK2O05klCwPA/LgDF+HIRMk2IC5wer5eSci
Ew3700pjCZIhO+WprEiDe7pfdaWIGMBqv18s/Vd1dUV1kipjj8olqOKVYBDEpmZoQm9mKGqqZbNN
ofbkmLQA2O9H/+PvJJDEMv3knTsHVMk+y5761xFf0vtQqP8t2I1S3I1pBfKt8Mu1F7T7b1P/nKz6
iYsGETKgDMIQMXb2Y1a/zhP15nvM1sE38DnPxX+Pj63B3KQUIfP5CTPFgBzdI5Vu50SONw92YnkX
WrjlR46jqHBdbyjpo0eXdnoNc205oZs9MjhAYENAw2A0FfnFsB2q2whx3NViFz09MJkdAllhJwZv
ebaywiiMuORcH3YLA7XjxX00djTDj2pKDecTh5zvs7YmPlz/s7HwECXKRLnQhLOYxc5ZZdQn3u9V
2KxeEyP3ZrZhzL1m/OHNHawDpGPz3sXJLTms909vB3JHDiVMuZF/VzQqgyU7/YFY5UhiLfVRQpUT
cSfU/TuE+5qdHpd9+BInNualMBL7SCV8pSXkYpLoz1lHDbs2ga3N3IuQmWYOkWgCrbZR422N6r0e
43LIZZZmBSMSaeMesluxRrfz3Wxbf6hDrqlV6/ZuI0X1dQCf0RZNDiMKug00FrC3fu5JWS+WIH5Y
sTi5a0QGaiowDjGmpoOPtoU2BwmC/EGtmcuCvT8Io+Fxt6BP0vYyNL8Wlw1S8HYeZxdpFFVVToYH
4xKdWqoN+oPD8JSspIp+bxNOyvDHwGdNGXfnXmOdLQgo6bLBbvIuM2wLcVb1sm4hJG4rRAYbCgxr
9wjuaWD+NrqGTtSKWL5ohpq7K+LozpyKIot5e8xeVhdNNsbRks7S4mI9q/V50zTruFidcVI3gGEE
cJ18XegA2YR/WgQAJ3oRB2uDuiHblCmWqy8uDyRIa1zWmmonHZgeiIY0zgWD5AVbPt4yoQyt0YKT
54B9e9w0oYx8o2krrAFvwpmSYfHqAJZyHfW3m3HSwkoqL1pJE/HvKfETBC1JAXkfW4AkaYAa3cJ6
2tmxbsqwmhVBWxx6PBRi+FcvyDXN9kH9X5QU3vdzCxB3eRBrgn11UvlK9GfVkEqtjOoLlNqD1sDi
qnZ8+OqwVXn7enY9zeR/kvzFXVaqweHTKGc7v4Pam8xiuud4d7nyJABKum0pjJiJQf80VH6r57rB
2qH4BNUJvf+RTlB9Nf4580TKm1B1oCwgL+Do1fTKNbyHPY64DJjRIx89EgarwsiO27/uz3eZPrli
VvdJ2XHtBeM6jlrE3oQ1DolEh6b+tczNfvOWxHjwrTIz5F5L6rk5IPU3Oceye/xgEFFanUJIYkkS
mgKaVBiRKW1Yx7/1s/380yBoixAeLQYomIlLgGZbI7U+6cxI/8qcelq38eS+eGKhEagwvRBgq34q
t0imAYOswMCvSm7YObNJrGOsmWdPRgp2sTzazjXDYXuhAKGnRnpDsoEaB1LtHAhhYmrAFh05BLpd
pLmcHOxM5AWKiIwEo+IUuStc8/okAfJGa3O+F6c/uacywGkvPwkEqrMDsBQlrUIaRfjOjwo+1g/y
MYM3izQnRPuo0dHx6rIoCNhx6mk8HGT8xw89VVcX04gKieB+hAw4gHJP0Cpf22BhmkBiMLT4a6gF
VcZnwAXnAFc8GIU3aec02ta3ja/gQP0NmsR7/28vERxlRvIWAOtxJ+ZqhK0WDXBbpSfYdz2dpl0E
kPAu5Zqc6NEAAry6SdwgdU0yJj1Wyg2TsQt2v6cMDA8V+QZ2x2g/LR/b2j8V6Db6kiMKCzPepF0M
w6KZuatMPB3tpdcV54YccHO+sX11Fy8T6DbIUEcfWl1daKoyYm5Amuv2sXDFkqvET5Z2klszaN24
i1XJFwO4FXMx61QcwvwoZ6jOoa/zmeAsG5ZI63Xl3furrupr8J7QvN/YQTEcsKH90kQcADBeAv4u
prIbncEtSzI2a30Pg97XKswaHC56wG2x3TE0Yhjkm/9VK3gEm5MuGRk2J3Ez72xNFlyLlkGG38CO
M/gnUjhh4NW2k5F8mLQhYdnuCelb7w26Cjvx3seXxc3ovqyS70x4DorPzcZ9u7oSTCgyimkHEowt
EAmbUQAhIsVBVc06AvOfk4RiieHda2DdYliHPA5erDO2w3UladD3TwSzovBgdLSSFWXYyF2uOcTf
v+PCVmGbFaogzNLKnz4zEt3D/8DSpHIAsOjpwSZLw5Cr+QA0lOYCyQkR49WDI/rsOZxii1H5bfyV
PRY8CfuoJuYZDKSLbjOKH31Q3UplqJ/2BnMyy/8PLyXGbgQ7YItR7sc4ed4kcn+2eNdGWOsdCgjU
W7xFcGp9VcgUlCGt1kRkIpIlZitZo7URgPSIP49ZMFwCsLfbxtJA9CbWESlMk60ILTQRgIwx3tzC
/XV6TVdSP6GbH0o0rKGzPGBOsir0TZusKgIzJuBUJrjCNGQhCE7gRP+wf8IugxHiLjDDYJuDFVeF
NsrcZWlFOrAmjUmbzpb08485FZmAT7ajLA8xtjK3rvKyM0NOjWHPbm1FvUzZFlSkVWW4EZEU4Gj0
SvWnZSx8kHTcr93Aa+O2ytEBz4ouOTkicoL6heTpVsmzGrYjcV792J84ZcTkmG3i2vmyzNJWsnnP
h8gH3IlqRnxS6iqGhQ8ElmhATPWRl+W7GO+0AnE6dLrY+HogVSU5FI4D0SqLilpTx5iyjIlui4ki
LLKtiWsKRAkBKXZJXKheRL07NGJc+20/1LBQ8NOndAWG+NpUy5KwaRob9iJNSohm/XeYVRYA0fBX
o4GIDiH6E64ZFjKKGemipORuWBcJyL69ueY4GX/jcL55CoAvOXbzla2nTyTRb1L/KtSOyP8ls7oF
sIZ+URTNkaAkvZiGn4nptBlFnqpz1BRh5fxIxzIvSVd3I0O9RNWa4TIckLQ4MIz/H6GyX9+iB3DR
UbxZ7iGN9sPybuK4F9GCXhpbZvAy5SkWJ4NIxdxgr1pMvbEiP56hbZAZsCk4qWV1BdZO2XZyKmIR
dbTrSVgMSNsUs3Gev3JUyUEwP/IslnjjK1Ncee5P9k0t4fDiBNKy4D38R/wUguYJ8fUgoE9dFC/G
+NBjuN8EdqK4x+dZhy+13Q5WYQ5b4iCJxVhexSnrchyZVtL5+BlY/AWeOY+yrY2Ri3lwKjkCrVIN
yC4Oxdkg4cMjXxBtug86siWkKmyDKDe3GzjEy7cQrivny02b7fLGCBs+XV0nI5doRlabYOXgMTw1
L/Nleuh8x4Ak0HkJVFQmZ+jWIwyJEIDWvli4XaUIjHy4tmiC4XakeJLv7VUGM1li8kGw5P9JIpU9
NlsZqBlGO9J71VKz7cZBaIe25TFHqEBBG17zeK6wwJR+Q208ZtNPw3Hz4ZRnORIrxkAcSAN6UBf8
ne6TnkxhUD0cUkmVy5cb4v6eEBET8GEIBcYkXzUDyEZKpsT8noMtdMDUsXnGB1neI4OyL01O8EZe
EqspSQ1aSWzm1iJTmH0sAh1t+qwBMkRIDqy7UHR7ATpTDpakNqcJbtrNPfOZ3mwaZoxcPKiGCtAC
bSl59AmtWkhIVfEwNtw0k0AGzUpDY8LSVrIfgJfi2tGybiD9z7919LU68pYDF1doSp4JxTM81deH
FImD+4RmJgRazs4lf6VGYMu3pBMRKE34l0Ym1azWPd7AHLIiwVMlly4B1rL7W0e594E+YEDQqnqW
C1Cy2pO8uEOlpwFjh9/oJlDv6OhksASsNd9mxacLIesBXHM8TqpZISeePhV5Bw2wN92hFHwGauil
PicDU+NX1YzwK7AR0JOvY4NcceiqIKtPHITzfndgsX+i8dCp86vcQpSjjO7gRi5JN83SuhPkuYcP
SUD++6HORj8TCEV2MSJSpezqSQ45WYdo9x3JwRJO1ymAD5dDVNkmxUs9IOHomuLFhStz2pJblXa/
4vOI87zL99SrYka08aP/bdS2yhcxouM2POiUGKywSEW16HhxRD0TmaP0uiIciVKxiRFWAhIt/ChB
oAbJatCOsG3fSeIP/mr1cK5VU4g7Te1LgzD/FsdSstghTB7lRrxZ17PiuS8TSsXSCq263/RoDU3c
mEB2CwjeLBoPhDk9yetHyQzLd087J76zeHR7c+6kO+TS4RdPPSryFieu48yb3JX7aEe2pas3QZOr
14m8D1GdMRBxm2KxAasxVMlQoOfLwD03GfBSBfcQKmwLkPbrEM2Yz2B1klTJaGTad5f9PzDI2LJM
aE45sodPfz5rVvlNsHPB4glkLyOHsqI55qyLdP8zI8zAr8YFagP6Wbj+XrnpmFP4+WylK5St+qc5
Nk+TOjvIY7gB+OmWRUr9aV41hsaOYWtqMU8V41hhD2gQQNBAJKGWiOJmI7y3DV1M4EiTEKBfl0+p
IRJ7R2R+23tdmc3q1quWdPyLWWN1/ayP8gxJxaOi4rSjbe7QXdvNcwOb+k4+BobBHXbQ7LjHeUPY
0l4FgOp0c9ocPzsjK2yz3ZhhJ5Pv4+7Bnj5wHsY7ETGSK8zX2v4XTeodi7CjQ3Nb8QoPqGL+rQjp
jmeUEjZiC9QlaGjmZd1H7WtYlPvsozOo39o9MCF//aDtoyPXaN6XYAcRo5vaj1EnLN4atKsWIrgw
Aw7XbwEEKl5uxeufiVfUR6dKlkW3VwBrssiv+2VBmvmDX19vAaablptcMt1gePsfJZWxviJdmyTv
/0l+cRHBFsQ6EzT5W7P68/Xib+zGgr70vTygcMgGWJ6j6F2cjjHgiFwEZsgpHG+M89DieD8sBoBO
B7kXNIWut4ez63KOtY9vwz+CaoQFdY8PyTDV2ASY/BtNEhNHTzEIBWVnOf5dJdPhznipHgbkNCfz
BSJLC8i30AbRGR6/bbgvkV95M/AQAzubpehOWUAc8SNQCQzCvGsEJP+2YhACgkr13Gs+WzCC+dtc
kM8V9z/CjQQWt5FhEeK4/qew1NGfzdbmABieibZ7F1N0+DMMzonLsrr7SFt6njAgGqdrF6j24DoD
VE6fv5ZVNDuOHILTxnsPqaG89nml2TwDMPThtQubTldwZB7Yb6vFnbV4/MPy+qvOcrFMdJDTxPBs
G3gY1Ms548E1ldfQErvc030DsNeoSzxpy1XYGWvpo0PVmkCjhI7xzNcQ03RtRv2c5gTrVUY5b3P5
CnwUmzSJ3vBlzsfTkaw1jB6Nrh3cxiHBitQvO/a3igCK3XUz2gF2V5hNMsF2jAHUjkqazwwX5Ck1
GB+xbsQLAAwHV8XJZUB0hM+1Yhry9hfc0dLH+zkHljYX/KZu0ok0MYBeDMfPvP0ThW964TyHH4DM
Dg0VBxuLvTXZBOYtPEwOBGtrIoMOo2wcwm63o3tmEecZcnOMgf4dksE6LG8MQDk6H11D8fYqYmrv
1E6AvNj27UUdKDpQhRhxoTav7pZYH6Ze/WUc81LhTWfb69I00k8V3JsqNugfoE7lvoWW7M+j3dqQ
+kNqqPI30O31Zy8UNxxP5WyWvRfJJSkWLq/ThdJ5J6CkAXVna4ADPOe3OIssZky89C8UCrNrKIrl
a+XyPbcwYBivP6vWY6LxYAuNSK9zCTpHS2KuE8L4E5YYdRLWa2e56429tWeVdgSDmxwxK0UBqsTI
6FIOJogdaECjbKZ7ln83D3lNUaPkl8IXDGAGdCMNhjchbmAvB9YV12OI2nhg/xLggZFunw3qi7EG
EIQdIvcU6HDIHEB+NZ4oUMcBiIeSJfzqAkLu/N4Xuh0WjXmbM+KRM1hdNiAXnb+w3W1qzYwjfSfA
aahBgNLc7lZMmNf/hqFAZIxyXg+ReMekWNfDCv/4qh3qABAqlnX0UYM+NpD/rXfdu3+P/PmJywG3
7L8GNzSV5WJ11GI37oDK1op4dJs8POaF2rAcHqf3TRY6hoRA+g8Kq0fx2HQ9MPI3zFnKdFe7Mlpv
uR2qxQLfBB6UZo+BObbE81pB847t6bAtTOLBlp3eojBx5OqqDTJu0qk9b+p5YtUKNw/gZAfS2Vw7
cBbf6qC+hIUNeqa72MBzbnSMteqZQNS+rp+J739v+Qacsj5X3r0fvxtCNT3ZDpoSS7ed0nk3POiC
PzK+/2BpGPr/6qh5Aj2WProo56mHpm3zN0rqN9Ql+H9UGGSOrqxwTFWgGqWN0syWV29MXEwgSdp9
FY5zWouFA1OmL+1OdBKO1QHIUZo/tYo6ByjP8RRO2CkYwBfTL24dVws5tymbMm7o7t5DHTQcIsPW
jFWeU5HwF6o3w0AfYPw0WfvrFvazVRBkouN6HCD901NfCShuDUbWX78/D61o1F9fTbl9YN/bdg8b
QdNgXXqd/aj3mOZqmLZX3sQyMhatcAUWMupglZhRMiWZ8otf6gBqO6L2RRHr6sC+e+TjwRiaPdoU
1NcYa1aVidLlHiqWGWHs5cR+bCXTyUv1Mbz3o2ZhJwrIyxAYt1R7xmXfV3aTz+zODTyZh3N/PPB+
kGcsyTYnz+iEIbIuBDE40UAjrNacCx6Fi3gox+Ip4YupH0j5jOnEWn5LN8RsgfUbA61Fq5VSgfl4
2gNTC/nAR8V10ctjM6As7gLb15HScduunUXCrGOyBtwKwThh3yYaVuR7zF5Z+p9trcOQQ5dkETEU
xCj8j6cMNaiYJCuU1vK0W9O9VHMLDH0N9lCXghqVRVJ0sJy9bXvMO6GwYi+HhcxC6o8wpsG3YwFX
Q9ucPO+dB1kK0W/ySBE7ZjXsn/ZKIJzUccAXLLuJ4x1b4TQiAlH4KAOi3By4OOEYVnixMyNEYJK2
to7YebcT+MO+TY48SuF6mfnfjU4YBV08mAqaEdeOREzZfTXMyRYGGUWAmwIehfqhb1oamLCfdngd
sTklnkyeX542JewL3QqZ5/hrnIbBvn+FvAz3nkPx4UtvL76QX6NO9vc/MWsS552YuNI/t+SzUKMy
KhHGpNkhqwT6CedKyw/NPr97UiPPaXGtdkcEGz6O4XtAheWGq6ETt54lJdD+avLdjSQF0uV/MqA2
/XcS8y96nvKk+sf65c7waGoinQmv++q6yRb8Yubql3I4gwuPBqfOf8CrvQTp1512/WOo/XjjUOi1
zPUi5uZpg8YVYH0bPD735DD/aPfBjmr6En99PUIVLOPMDr0Rk4cPoa6GjYwRtL2q2VjxICQgdZc2
X6P/9aAr44gSCvYKTJ7l09fjUM0+7It7coNKMI8TnIaUGAgmRPnh8p7Qtyt4IK6m/J1FWo6JyWeW
lESF+DZsK+rOUasiLb8OII0wf0ah/rnThzv7LyWVGLmtbhLNArZt9A6O7w//9gHxDFWNTG8wUKgw
DWSpVFtOABdMxHFMl8f+zmPEAk3cQqJLaO15AU5F1gqrbEdmim/m4OiX1Mf6jecNk1wJVcJSImqa
vuzchQMpwrFNJwYpBKgZBWw8/UkuBOiOmo6pEbhNPxqF1QPSs04VUh9Q51y+LRfdG2Nuu1WzDQb0
vf92T1AGOKOrkcDXig4AOfFVjX+ysU2d4ZhNqrXUDrdbbt3iv7jsKACYazO/cPzzh12331Uf10jH
VdlsMASgmpMtLCSdv4GITmYw7+9cir5aqVjM4eEklnsoshJ/iKkrfLMUuSttNJSHUnt5J5MBiDrZ
cR5rdaK1r8wmJZDZVBqOUw/iZ139edanfPoBHW4DimUVeiH2A5mJIfNSOZo3DQRmdwnwG5Db0Upt
N+bQ4YdgsbwAi8Q1ASph2PVv1hXhfxrPv6UECvEaKeSyH4i/veadS125uLem/gAX6VFcBWObHc2Q
owhVRl6FDz7v/9h1OzPF57khJyKdbjncm5cSBHVCygz+q5Yn1sFqP2BvF9DLs/t6ce77bk+MTDsV
jrIAEX/uV35mhES6xXdZkbgEiwD3ojT9AkY/EmzpFHvebihxo77f5QNO5ub/7KCh9uPavmeAl/V6
F7443Wme7EnmJg/R8lC+q94Yi3wFzDq3tPEG9qpJpad46zzPxN2sl7533+DRtKU1BgPMwV8FNQI+
CWIeGfPGNWjRzv+f9seVJdbABZDADz8GqRS91o/GgAinY61lOFMowjvhNclhjYkilLWr+S8G2gBA
JomNwjn1xCdyvHaYIJE+O1M77z/d7HEdiEpc2jJ33RyoMasLUYuIfln6PWP7D2WIPxNsg6BkxNvY
d+6YlI3Z+h2GoKDtiODLIev+vF8JvqdKX/Ast/KG3kLpiayjH2P42HonztEEbqssdgOSPfLtKXoG
nDQVqyKReehDsfVe0I7ap28Bqho2PwYFJH4pxavmyedCNjav3ypULELGkOdVZuNpZeD9sxhKONP0
n5tnYllxIX3irPd70PiOtCtoAZ5Ix08U1IOMD91Y2dljTbtm8fTZUtpS8jvbm4BQmA+9jRfASEbJ
AZ2kZQBL66zabRiCS3IZmq9+MQhoHPjdjuWzUNx+28FZFJGc9c2lwp9jvna4vfzDbEhZSKcmc+ZM
r4BykCZard8brYp++iw3e1UUacfXG8vZDerD6jFsJQzPpqeyKzL7VFSlKuspS8gir8XmVqpkNdWi
uNhTMpCwoUDioUmzNW53uD2HWx9AzwFNN4K1s90gFUrpyJmnfGqocnUlRXn/Gc1eNCrKZtfWWcSS
DZuQeeY8COAMkjO8Itpnl+n5sVcRHbgmuMBLEJWfRK5zqoISVlzNZ+K80wHOuCvS8jTzxgsuvcrO
0rljKD1qVBkRPmercVvyhhtsy9a6VYcxDAq5ojyw8nRkq5WOSAYvDedWPKn1GKF8YnzAj1zRrDBU
vvsJAqT7nGQ2ZKx3+re0YmVDyb2UryZP0xgcuG9tPj+9o5ytU3aQ4hyTEY19BPKuh97FM/ZzQYIa
YPc0lrTztoJ/R3ozyEBc9LMSSeoaBa4ihZ5atNkJp45CHynKzamaVN+Ooc1gLJT5j+nNgQf3lP7t
n76BFr0Tgx14KryMx+EvFi/x9UvTjhY6Pz5wr2rHnftnrKKXm0U+jhtj3UIfiYPGlh/CNm4MRVB9
VlHSUBczcckFLLkpasLfhnOXGrFhsytQ21muZ/srBJGnVSgIodvttEkHqmLAOdfBKfZkjswuysEl
ua/3wkxTeRT2NXvbMzPXYkdmANZHjaTw+XWE+I3ClsqJspzHMLpT470YUjVJCSEanUzmHnWKdb9M
J/KMs0r/+JXO+2kTetVt0z95uO8T3M6VhBU7vDuXuOs6i3bpCmgFL4MY3Xeavv8h0U5RtyCDPsVz
tXDKrlzD+RFCxowJFpfNC1eDGZCaB4hxjEhLy7CDr0p6OOwC4C5xBIHvn+RafmlwiEmeBr2RhhKm
wsJSUr/8eCGHiKGgccSuFVbasddaCjbbPvOUI0Zj1pi5UsgFE2a0IBDLVz8UGFXtxeR2gpTxdV3f
zjM6yvYUT3qsoZmwRDfxm0GY5B/0/LWfoByyCP/FXzcKwQ0E9Lu9UQF3Yq5JZBDWM/50IF5xAXvB
GRbMyPnEBmz/cr9hPek7dl9nduJSirClIWeyoMF+ol/Q3ImH7S7mKtBV1oKJmGxNT+JKaNInWNef
3ExUjYbFywXqpNsX3Rv0VQCLOvbKh9dIc8BG3+BS8HGSePttVaa/RXabxSSu5Vosk36Rrsw33Z7r
rz40KaNnUB5LCA5Lnl7P6wZ+TKzj0slQuvroMTXl4ekr3CL1s/LGQwWMW6bgCPmQXWsZ7nXeoIXk
eanrUn2+srwYXItNdz0qQBDP30U5TzQAXN0wS2BwR3VrPVHjOKXnVu4r4HqPku5THwKKRjfKi9p5
t7D4xE0Ndy/34HfU2Zk+oqiOYn6ZntorZGrxQxVZASRzRGuwmVq7UlfCxN7Hsg0OezWbDvnyIdn6
CLRDSSA3Vf4Xz2ReiBYxZ//2l9AlV1AUxwFFYGKxcflBB55hQ6hEulgV3lSKi17SsQXUzK4ibpc3
NyIUuavrHvd2QpAKGSTfkrdMh8hhmukJUHznFtMrUa3W1+Q94LVwtA6zkL5LW8F/oTFfTkQRsWht
c9Gqww8zGIWt681+kETOEg0oHSzhsX8JJLdsqLZeWMymt7W0GVUR++F7CZfI9ouGVjdkG/ielkwt
dZfYe+iMMp3S4hHly8xQdHzSSlbiXaswpB4v6Wh8h31TJ6cib2biVu6wSQTLqqpAlbClIQaSk2iq
wQv9DeL3j7XguBgRHiWqX+wox7hxR98+0ZhpsU2WWv3qlEPbdOeC4EL7hdILCn6Cj1grBw8hvazI
ozejXX+3mRTvLZFK8mNnkikOO3V80P3J4HaH+QVrn9P+Vu74I8YDR8IrdMF0QnzjTsW0VdupzTqt
hDy3Wf9evUO2B8YVwX6waMxow8d2HKxWeEF2/HnjvWNGyZ2iw6z5YW1dvjOPTZB5p/gCsLJluP5T
gfL6pirHk7nSuB4vGR0W7vWcVBXvJjk7+cXYomoRF7gCpbvZ9T0e/Oc37pjQBNQDGApQCtN+cjp+
5TGY2M6V8pYLtBuvQxI9zOWrNlOA6oYKtfyrmqqiOkw4935gJxYUWJsTRWFJ5bB87ZUNc88KsUCn
wEvYsYMD4TFp1ajd81tf1U6uGT3l+ez4V+z9GjtLoIFqK5l9OdHrb6vJHXIXv8RBs0sg4D61P1Z8
7ZsB2l92Eui8yG2S6hwpkNSSMkIcJIzImBvVeQOaoKwsG5gOPgmNQBuHkKb0+Y3oklRg7EQyzCtp
dwhOXceXNkH8bRwFHZtUMUeODf47QETnbfHKDEG4erZZ9mWjnEtmvw1U0MwHSsNjfwukbJQmdeeS
6zW+LXSscYO/oS22MowTdK68yB0/RhUXc4KAf370mdOgZ/XSnOTM3yTUBMq6L0AUp6ofT8uiYYHT
tZvISeD6fbnV17xtjYwxSP0z2Yric5gSB+XOCZXvdKQMPaiLVXrg56Eu9iPXzeAM1nzcbnvT66DP
BN9Tvq5/8hX9MO1feGtB7vIV6sjiptRkjPqsbEB74M3Eh6o1qQgB1oncoXVCca4DWugivdS97wlM
Z1HYSWKynedXoFLBuyuNp2J2cE3ilPaBv+z9r420ZBqhd7ojBRe9U4fPMInkKEJkacTnvbPi5wpQ
14ZOGLa9AEkco9ncc77xhOD/WluB8eKYjBKl5WVcB4L3CRkY8QTWK87IiOqCrBur01Y6M5fPwXCD
Am82GZ2Idm08UhPjz07vSULbzpf5XQHkQUjt2I07w3HSFzowUufC0AtcZqF3lqrxwndqbJVyCao3
JwbdWd4+VaSxn17wCpu3Im2WyMfsPPWaUKSUj7PKLeTR6NRgkeI1RrN2bRZbTLTsBADNle/eu0jG
YEB0clr82X5+MZOOmBexEow+WQ71XGxSgKpiheEkRa5Y2So1YY14QnKgf6N2iX93/rHlaNBorj8i
5jHzBwZAeFL58VFyJObxBQUc06Y6iiByQ1f2mDsunp4EQ2IY3hYaQ8/2s8JDjvHITe63IvPKuftj
PXwmvlmHmbmoVJO4PC0AJxkR4dag3b6bEK7S6+j6Zm8299DJC6YN5wX42XIMuN/3f0rCmp00Ytji
ZaEoktHRNG8rBQxboW5hJqX6sMUCiFsfDN7YB4mdGE7t3hGJwaUGvfEAfra5GBIhAijjt1ftPNQ+
ZxReXiXQZsOsD3w8uqCb4ItUhYhMboAbtdIerd+igXIk9F6eaJp5QjVGAUAQ1KbK//rh4iciSoC5
3LUUJBTGJILoy2TzKfHRXhisLKkBxsBig/6K4Iwq9R1UbC58izfnZ41zVuhRiS6xZCHwYbVWghzb
l1PvI02A2jLhCijgeQydJJdnrnU5ZapZWzQa7LsxfoASLGhjdVDezz5C77TBarNV+fcK4xTxYfOV
g2PGlFm1kq2/8KCtBlD+kV5qQGDF44XLqxGoCO+NMKAoLxqHf/t0+jWHMc5x1/TglH9WPZ5eGQaR
tDMaztHfBAtmJgy22xsf1h6P9d1hbU23m2e7TOBd8AsUWN4gkFEi+11Fjp4+RHUF509N93IyCY6x
qAJsLXUpgTy0nixJShklgBlrSYemcApJbBDewtlbYFqxaRtts8z1vZxQIvmu4S20LL8fLl20Ve9n
RtWRooiIkYSnSdjqCzfE2usPz4gS/5tErlMfuTClbNQIKBEZHODtR8P7jma5t253ZZwWdKvy4vmx
VhphzetC+pLahT13QUplB9DJ/SMFLh51gk1JQAYWIYimzdqNcINyIgwAjZaY8GVScSn4eSSdxoMy
Ja4BUvNema8R9tKqZFGrNHHilANGRxh7SFMNOyoyIY6Vr1s+WkS7D2fKrzDglV+y0s0uFPwwWaiH
CVZRPOUwtmZo71j17jU3asYMNXLNis7dRUq2I353y9SqN/P9Z6vS04X2IpjhqnVh4RtjVBcrkB69
1oy0OyX0MS6bQa1edQ4zVBkObUWWsScho7hmWBLl9q57ouGD9KRObE5PuleHgUJLubGU1UHvFkYi
pIxF5+PTHojbQ+nTduAO51xFAs92g7O+ZixTTzncAG/ytW6CozVnMBnegNL/nTGiWhuCvVcOC9Wk
GyBGHq2gp/uc8tT9Y1+Uhcy8MIqfBxnZn1xNs5XfbViytdlI8aF4JGPBc4QXOCw1xGKgG+LF7TT5
UTCtD4Ep/gB4/hQSWE5m53lDiJeACTQW2NMTKJ9feqR4vg0b+eKu1Xezjsxs+CPt/Z3/0V1h8i23
ir1dqydYKthyOGKr7qZhg1mO6l7A95F+IBlvBSXKq4jrOlTsWbSDJ+afxLQd9mBqsM1XmQ8vFxPn
ONT5AJszUEM38BLiJprp5PEgVhDuJWV4ovaA3fXMtsP8heFOvFvXVLAOSOgBlAadjjk0v9AKkkMj
lpb0F+l66ZdrNvdw3C3ztS75KNwfL43KLUyb+6e4mSvgFz+W65eV66ASfSGFWZT4S9aTdI/GRRrk
Xy88+A0wE284jmKV54H+hY0UmEx/szdMsnMAdYt6ExyN78q/R/BDW9UVc+wGYO4DL1DbG26feclQ
h1OncGFCSa2Ftsls/8L8QFyPqkZf+l852yU1Wms7L3iUXkbQgp8I0kQCkIIyHyCC9o58VtbZyHxs
tpil0SxFMXBRKht3+Cty1dBrvsvRPPZhlVyy9h939D8oadS4NCuwztAzo2DhOFeQT7Uj2DPpIMeh
sfN5P78dB78eufAci1Ff1RAnXRLXnZAvvDsVn4f5l6nBxuBeCZNrsKHWU1TiKmcfNWn7/m5vp0bw
B6uQo25Gn+0NvHT02F/ALkThSbvu9vLdWq5hUbM7mbTM0Ah0fGHDeO5FigpKEDPBc6+B/nWxUZcv
rGnq9O620rrofiaTSfD4C9AQLk8201qOICtU0KRfqJe+hKdY/ss0O4b5BPirv6YiFUG3WR+gUSai
ElD2VJWzldv2yeNlvK2px1T5RMs9EbkT4XvaxVU04t4AdXt9KXA/flALQy7ZeSOQBz9kZvByjSc4
6nXndbLDjIRY5qUu/LHLz4O587U2vFWDe3LmUSnZ/bvGW/rU4tWDuML9trJYk+1iy5+TmyQp6qQe
GCn9I3ii9HG3q2hmooUxjSwk0RcKkUbw9XZsufNJ4gzOmyox43HEJxcidZDzIC7A9g92hQeMbxjA
jzRD0m+MqahjhA33ME2NlaKpshlYS4qBIIb/5nFcNkDAoq2JtYPrabNYLNKPae4ojM6LTbPn/aOQ
+3+yHQRZ4imU/bZfDD9cliMxgdUhYkoC6rGnM/D4d/oQLZKizC3PrEg6LlxmsMb7q4Sx3oj6oS6P
T41fxFyN98HzgmxQR/wyUDrNqLUnSTu+1rjyx+Vja6dd117Dgc/utlYcdRkRauN5zxBaRJpOm1mn
ztKv7Uq6B5y4qMO3d+qfI5tP7rIgbllxHxWXPohdyhcwNTIawOjUsYPd/vefUpm6FySGR9nKeIAI
tYewDYUr6za7gi/WWWWTZyVCFDQcxIwDLpz+MuneehHIeBTDlvNTRoa2DyqEJRvpFpPYahzBZbeb
lc6ScHXwjL5asILUvO5ODrP/uXfFOuoli2D6PlrVybWOfPkUBECDl6vfFmBE6Orz60DuXT+OsGJV
f66DrZmCX76omrTV+SdMQmYNRqzRfsTopDmkMVRjAQThr1ISxoWrsQSirnL88xfd2AWwzBMlK4qB
9S+W8v7EX/QN7drztZBuwPewUXBEM9T6G3YPMp8k/Q0hIfuc3EGK7+tnIs+lRNwyMMSRbPXa5rOj
pOEifn4OdFgMt6ybEAQw+4HcIlDH8RyFBaV7T/apNjVo5lx85zZWwfmTvQWd1ICnIk3/+4zllor7
xA4aVAdkuXh+FQSfZ8OkTHihfK53iijquz4tcqAK+AqFUB7KxIqje9Bm6EquNrQ/0jJ5OX0m8dW+
4Tl4ODykj/SpYaQwK1WofSK31S3gVAxIIJf/OilWgmhTUCtWOGizzOVfBZQrkyRa7Zgm6w0wthsp
d5V92jQSFQmxHJUmvK1ApeNvQUn6iNpaWO8a05LxsJ6EPVFPjPxyttpIkeoPGxIy2rwDlGm+M5C7
NxmeHvESgyIznW7xa7fYUVUdvDxapJBJVTGhuRlPjjPkayDlqFoNqQf0y4Dq2ZDWYKO8TDjmLIFz
zTKSNjsMMC8Urxg9LKGXAPVoukQXBb0X0BDmR2LxJS2Y00O1zSauxBaYM65fEgWqvWVdEnw/HTUv
6OMdTJt2H1ApiZfPUkFGpBfUGFAmCjdp3UY/MZmo8XZgDiw8xGDiZeN7F2oENBeWDRTkZhP7edkf
TAErm0Bpn7uBJ7WcQZEKec7VAbMVp8eso5yPgit+UiwXYvZBNBjgbiB5w2WLOFGNftMpMlu3nWOL
nmbnH5AE3+Etwqcr87cVtp02rzznyvq6kRh+VQmYz/6BufwarW18eJUs0pa8Kzyhl6q/n5z5EgCz
cxNjZeBXnY2IKCcUGy/QILj1Niu6SPtQ3sWZzdDP+u/H9RADCK19D46TEZjzzGk/fSwLw7oeEaWm
I0ZtHPC0KOUN/Tz8P+ZXngPipdDOfxY8CCAUCYe67xpqa98DMXC7sCylB2AIc6RJiyZWQnHjBO+U
zE8KBx2G9HrFTzaNcqJBiDNNaaiDacOt2lG377f8B774NmfQrrob8XhEv9TiYZzk2+97IOsikC4F
oz9O5fVz115VNCfspi6b+caMpGzrnuNHYnUhSV702z5wbdhfpdm+bW59iQZEgRLz34IrxD/bAwTt
MpSd95O2MxQ31+IvPdogUY1GK3jhp0Oa4hYHZSy6d77e78WCUvL7BMCyRj6laQfamWv1re4ApQ9n
vDjx57BaD21minorldKoPi06Heiz1WFQA9NTaJobtdToiQ2lwjXYcMBn5Qd9sEgcVSRPsC/6LofC
lGDAYc1RHC6QS8bQG7u6hNOKq8V84iSbs0ekgCitVAH8Hd4pmhqCmHxO7WdWqq1aDTC3Qqkx6nb8
rgCqdV5wuRvDOv9ZxPBqS8FzXnCqYJ9OGLXRr+02zMI4w5c2noGVXeSkdp0ACy8tDGw884xJ26eV
mrmsxjI9HGl3r0+u3e59G0DfApL8L+xuqomwgtvDtpidPzD7PP/0tLsX5GheypLS2NbCdnt6nyDn
kwaO3xa2goIh/BiXg7wy/cezwxNEubmfMPCsF/isQLO7rXxZm0TiHdYE97nWZzUTMy7f4KCJBKwm
q+cNRPgtq/sfHsqgmYp/UCeDE8DEQAg+F+AlL4x+91OxXWnScOH6VILouYvhBZPoHNGWb5qJEo98
QQigkfrrKKrNfsP0kCI7eXaBoWW21jOAfLFlFWxjoZnGcyqZScbUORWDYsM4HfdxeoIEZqqoSulI
DV5snHfsI70478ktnnZAWtyL4lt2OLl0H507sR3ojc1Ccr+hWJv8fW3I1tb4ja3IIyva7SEFYz/r
RLuNXbgzaktxWb1lQT8JLVIy2XN24eBESsf2PbB6hz81zoTssBsjPSEopZs0wW+fhDDPTZWUwG3N
yIVouw+zl1y5w+20uMfsVa9anobuZSYKfKxis881Nq0NBtkP+iSDJ/IPNuJfo8R5oCGzvfnGFl2p
myUeU7TdGxraKrHoXwttMNAqMCGxnEy8gSX6h7kK0kcrMQU/P56W9ENPJ60dCheH+vcDbc5CbjHf
rehqwwTS+u6wOdbqmJxS7Zq/C3Fx5p0+umM1U24ozIWk1oZuXgX5SCJymxDNrriOPWzM/bPBNg67
Qu9yBSNO/DgKrV+hjUxqZQ2G8LwSTCORg8LRVTeabNha3X+eKzC3sEu++f3zV/v2rLhg9f0aYXZf
+ma2gj4MrKtTxwm2V8x+ZHe8jRFuMJvVxV9rQ6iQZmf2K58mvUeTCWLeKlPlCj/8CFvX2LF9pvA6
hEI6ZfQgODGbcUYI5Y/JvvuDtxgIUJzN9xi3dk8Ui8No8BTGxOt6XlWJl2PJIAzqk45UR1RQzeWw
IUXLtUp6JA/sNIQkngUSh1LBmdmRJGgqrPz7IUl09DiXCZ0NxmrHZVAZ3gquuSUCzaDx6WUwZNIU
hAF1E6blTgOG82lUxLx5PFgzl+tBgCWHftudiQIMJIFga1tHO0OajlD4OCnXQvEiZ6wSNzfyxua6
WblIGCH1Zank3RwPjp5UcqI4S6WuEapVR7Ps5rz0bebwX33G/S/mAABaZy8g4Dxc14AUD3LtBeio
MLP0ISNFlKyQpTITaiZS7xKdvoMEetyG6piPTZlV4HU2BoLTz9pvaswhrQDgfFvDy0V3nplWsRcA
JeP1Yroe6N7Pr304iHZ9JY2E6bQVsY3y3No/8m3YXw71DK5yMJiuuxe77BjmsWUWDk8yzGP9A73d
VrwMnmgTcJCtrKay3ic2K+74KvnL00NkRNIWSTPOqiynAkfbXcFmGj4k/Oqrvy+TQwjUMk9F04We
zT54WrIcSajB7agdx96qIZ/YwwtnbjMxzUHS1LGxokTFXXbLH01y54EpL1P4C4Z5RMY5lXjBLaJR
M4QG2GNf06PH+2nVsgAPwN9gByAfqfqnV4t1AGjuIddJwMPZlit0U92pk1bwVBxRq9SggAaNcQVo
V0G0e3JakE+50NKLI5sJjGnjwQYmM7rg3Jkdq+n8rY7aPl4y4/DIwLTv3v8SaHvRaZZkhDpz/q+f
5zRf613jopU4W/V7gtf6J625OFgrh7xT+0mU96pj5ZUFOj9d1NU+6u85raJlcbu5iPdTfM3kE6PH
cXs79hbsX2U2GMVe7reD8Crf2Rau7TyTO7Sspoa7iBFxKFzu6CIFMWiW3lB+PLB3ipGYtlitQ4Dz
QnrusRQCekMV0QZSbCQDuuQuBCftL9Q50DOnNJLocau4HseKbkt6O2f4xTcmlJ2gpq/JzENSnR3b
hyEI7/Nh5LIhieMGXiOyGchnjVZDxOIbbOv/ESBa9VaTsWcG2fmF55D7zHe3vg6w0haSmEJnau5R
cBCfsVuQEdDvTi234RJrtIzNQSAzYlAjgaU5+yjx145BoNaX2qSEfxEJIzDeR2jkO7jfht8I8eyh
zwlJK/kUC2E7kQ0j6b7WDKFiKj7vIDhhgyF0s2dvXlb9cfnaZ4Ok4SLaIW2RDp09u0T5ES9CnKCv
nlTs+LfT8gEBZ27xMvHEb57tf3bZOaM6kK0GAqKxEeLV+gRaFppBrtyPTvzkXZR2PhW4d39NMvuW
I01wv7RB4zq60rWmLUBXoQL+VA/QnfPxXbfb7py5TnpWljHlcAMvZesjseLk8RUOTvlPzovBmScz
lhwE4Ga9RNZ+RThSdcMxDgcj4t3MPXjMaNppIVYGvCNvT8/c3fZee7IhdRG+Kh50mM3HfFnZEo0j
HioRA6QnZGf462ukImaa0KJ4mZb5IHcDL5xrDgyn2jOrZvOqrjUlZdiTXr+c13gal1HrDzVHF7yN
/GgirQTAe9CYy66aAQel7Ha/O/70E8Sw6kZX25QJivQ+Yp+qkqmLRTNYdjaB8bp5F/murk8FYaPH
gvYuUjP0vfZ+V3223STDso1BcXRv8hblRVCdeC/SOZ4V5zePYfi8M5RkoP3t5XixgT1puh2mhD2W
U8VN/hqMEDM6Kg6NMqotqKmpuu6V3riDtDp5vWPQBrecTpSfD3ngBlRM2EatMi7jTxndTanXH3jE
p3w4Sa2YedqT5NNJmD8DUXW/XRfHXS5BW/zACFcjQK/nJYTXqxcM5HT8KxpWGQajLbxs8bgDC9bj
VA1x5BxhNK7juc0Psep6yFjUimiF2rtDTvxtPrkMjoffKTM2kQOx5CDJbxMR47G3QD9KsPMVaSfG
pzh3aKqT4TWryOQWgl74CCWnjQ7y3MYPJIgWw7cXxT2jW/4w2hiuU7WHKqsLTgBK1aMNzxkQj/pz
5W46fLdtFnqm8+++L4O2+StHwY848s+ZKiONLStILYVvYR+c5AqJgSl1RfC1CmoIvuo2jAfvqlZg
N2Dc8tdHAN3qp8fUi4LQWgTz+A+ELNNQM4eC4Q5ixeiVbhABJehiYSsAb0mVP61YVbOgqKAv+OVG
EIwgneUda+ze3SO5BpvrgJd59ewD1Qxj6lQNjpaP5Ma9hOX2fdnhEgQNBqSqPGBnt2YqixoxweIg
XP3uEWj1Ig9ldE0Csd18wPBmsMBQVW8+0LnZFK+TmJFLpPRYGo61xJNn7PEY2me2Wv7kDBH9EvPb
iPSxf26/zFLY4lzJp2oRPcVgCHTtqSGYkx0D0so8D+QLrXDpNNTEMH7VhDKitV6+RfS/C941RtTM
0s42QZkLxv7+qrZ697e1npS3cOUNL6rOiYAM59TivWUPmH+NpNYgJCstiexTbzwtfyykaEAkzurC
13pwnstxiszAYWEZ7jgLIjEXLUHwnRpXLbOyWm46RWR1QQwyWRIu/U2Chh4tJT4B6SgsWqq6ciTN
MZldqmSdw6Zr7S/LSmt/1TU0w4c+Vr8BtgyVnz+qggY9Ky0oAzjjok8JWYBPWgLR1WowlMigFruh
wUc9UDabEvexhQhNbVmXZZw48uP3Iex+js71HcKZbweWQ1o0Dp0x8V8omcC8YY9BSx081Gnkb02U
opNu16EkQ+cnTkxqRHtodv5jx6TBAD1oEaJ/EbEDM959WLTKvc8hL23nGRONKAIcgCQRh1pOsiIk
KN4P4jyxy24jRhiuTF8CSM7ewKsxqU+fqq+r7Ov5pyjMpt5zo8otpv1ZuQkIrTBm/Z5LJ+WTnSAj
nB8k+CLLHHUNGpBg7Z5obe16+E6cqedw4ecXDP1v6XhkGzcpO5w+Bxbp68Pj/dYkCHcAGKzaqC+N
nCAEcynwyeWl6+mottxVzaOsl+jhcWUAVqiERreq0aZGUqipqg3Pcwv8PkXpSgmbtY124tjsGgf2
Nh+UytwWre7cUPzIS6jX1+CP0offlRxpwGjUAEPtzMr9LWMEtdcX3O1Z4OZfk/uYiqhlUxQqZMPN
2Vr9JaxwxC+S5Wf47umLvNEMqLMGX0vPOi7UkKL4PZZ6IUu6vwT3lbESqO+a7IoTyEH1rinn8Ffy
DVNYwWib9aE6Rzvhr9XetQ70gRtY0lpdZVxTSyVegdy+Sv4wwIq7MXUs2AMeNgaCRSIrgGXEv8Ff
sfdON/xnIKvvxHqZcOpSyVBfdfovR5mdNB8a64h6K9DkUvXpEiXJRKUSDsVpXiz+A+/9Gh/Cdru8
rSRDTiKZqeOkYe4OCDmgF3DQ8qWwC/9OXOY8MCmTBb1epPn7llpdvvRWi/cRxMjT1NGf6fbAptY1
qjBUZb44dJh9mFzSMFFQeItGLt0xSIf3cqD9LYDNo0I/qUD9VgzlqFZ05TwA49pszF3WIABYrkUG
Tta6xcshSxiVrcRnQXzF1txE/rjujyaYl8B3yUNR3T+ue6HMmmjIBvL8lyrRpTPZ2AUvt0NTDpo1
LJ7QV98WN6y8aIOXjvsBHrvBqA0PcVXLaikzPDUUR4X2fhENTp1CP03JKhcjqNb3ZrWsJc10qg+C
7rzS9IKtwiRH/iW6+8PhNpwUo0HUV2wacBO38ig06mrQcFJ8IVQl1Kat2YOxrcftQH1bO5BGJ/HQ
dh7IZUTL7+nXp9x3UhIf2Xvxeeafju9wd1280EqJSqVSVvc6EJXL3dT9wpeZzz8vOC02DXGUxlz9
W127hM4vSQj1WrtibAUDNwxaTViZmrkywUz05/d5+WQEbTQRGh8ViZ+tsNv/Z+u3QlhZaNcNw9Ij
IXh2hLg33Ixy6fguedRrrZ5XuPZseekdDvAe2iA0d8wXTmntQoigqlhbChEviTgPpRa/Ra/UuJ+w
fGxPsdnSj6+Ym9WDNmMsRVqpMcZWijUl1RshPpkTDKEDCvAYTXNsDOF0pT1G2Maa4uT5kQFSh4bP
z8999Pt3mnA/4NYX47PY3s9rWhFqLnyxyuKO5gxFj3RdGJhUy24lvcO3HpUb/lCjHBa6vvOgFrfs
Zltxp/QYCPtBcyk5Qk5rGZGopiare6UAplobpDg75dGZLv65MF1M09/TrsmqJHv6/LgLHQSvOkjv
cG6d/xhZmeFAZu7SM+U+dbl2GYw4PM33SwS+H5rOWhIMv10q/+cJFoAzzIxKK7J4+CExbrVMdVUg
yUeqrHecGoM67Viyf7g1mUa0G7S0KWhhV4n/qN12FMCkdOJF8cWDiynB7NBdIjuaXXY/rEeZ1434
1N3pkvSoefQnQbwuV3kRsilz/y02z9NXSsIugg1gMDFh1hn3J08i84wR1br+FHZC0W0s6/wzOJlo
/gBcpXE7NZ18n/hzZOhKmaXxrolraNbAu3W+Za8/9pHuOTpX8VXuUPVArWrnVvmHsvF9z6wcGlXj
GGc18Xm5Mraiclos2I6q66AI1lMFsnYSlt3T0zT/p4bSBBlgP/RjKjf4sdzvDjb6uS7PSLWqK1eh
OSf6/A2uftMJw/O+wv+QUioqRckzU0Zmo0HN5JaYEDLZWFnflQFg2kce4Lb5kbDK839/5v8LK91X
A4JTbLlv7CArXIcT0I+be50BoBrMjvWJ/ZUeR/kaVoXGYBAIaVpE/frqfj69IDh2a7lRC5l+VT84
fnn/U0ARL7lGa5RQ7oVOnTiMeojgcohpyRvDe+h8fBWpUwqye617rnAQsvn2vuA1YSkwAz8Vz7so
4BTmbEMsCDWe66p77K/YZq8fIhe7fve1mncvi4wbBJBhxFTb370su45yl+LdzaKPWJKTuBd8SLbZ
GwqqjxYYytlhm/tycHRB2RB1zVK6YIvzvO7BXfyZgAkgzQRtPVlyxiZy8Wu5Z9vGEGk+hYIt9cLM
VaCY2/X0fZa9jbkKZIopYO/vRE9q1/sb3EDlMWOXbDlQUaBciw3Qgv5fG//z47PCZbGGgL62UlHQ
IWDfm39bRWQMqFJa3z3lwFi6M1+Iz08QZUS7nK88SEAsYpdB/aIG41NB9Ce3mdP7azTH8PJ0gjHC
rY9nV/8S1fMp2Z9Zg+pzaRJ+ps+XKNZIFwoN0Pl7WgoA8ufnRnGFEP0Nz0Ci9Gf/ReGiKq8dD4SV
9Alcqd8jmIH7wY659K95u+2aUTZqlZsD+lTHsw+f9yFCV04B7xlDXjsuPpfGvYxLoJUwianrAt+u
ChmbG0XBJcbZwKiXlwGkv2RU4b08aoxu7XWTf1nFVEMbL+10gOty4Frqd2+fiNmfhzDjjpMNHzsu
WVNJ4VISDFxCzS/MVdrZu0hE5dcqBC/0++jmQLEGbs80l4GJMv24YMwyXjTWBileuw7H6QdF+bOU
fo93oDKDTtiqWG2De3fvghM6iosmiAu9dFuIpTK2qK3eJM82zZ4arNTUdbO62ws7zJI1Y+v0LBS7
2IyTz+FEnm+8clX8LENwd//yoC66UvIldglnqf+ZQdp5CiUH5rLtSGkjC0gnpBo6lAXiKrxdGm1A
XPvTSIOZdoVj06u8ic3XC/et42LjpXcHv69OpIM7tYyqLRH4FyaMMgu0JvAgfxnlXGxbz8EjaTGc
jlYWdTkdMaB3M0z1qsS8gyRL3m1mzV/+GblP3nnc1z6x9QSxqqs/ndPOJQUNQhOQLARhHt0MRYgu
rZ/7dbtQeLgXP6+eaVUlEKpjaDxyNT3kCSK2NVye/eXTEGtZd5sKFGpYHV9XDjba52DLzdUonFRH
PzZD9UL8+hD/aiItjZ/x5/zM0LWA2Iz5bMZ1Iwkdwm1KWlF3SPBe6CgXGGQ4uNAOdPjex9IlFYCt
wLWIUWlWNNqwutxl2WLG3ZK/DXvEBigSVNKAlASMBio3zQVMjzs5Bq6U593q5vWNjIhy1pbqzbsQ
zAoS2XAYJjHbyCSVeqNPEDU8JveoMzLkL9ycoIsB0SKaGlt6FIRbbhUyYIp4HjPZXpHQ3VPgyfXh
PDfLZOnHYnIXgxYsFZByf6jqRGqb3HbW5akNYcO2SvD5wewSkc+8Sbth6FyHZLPwu8t/LrF8kmYn
crk9foLWnEebJ435JbiZVxXYygUXAr6ms11RVgBKxzT+l5uj79vTXoDAktaE9Q3u9WMEG9xyffJI
uh+H+yKGm2HOzdi2dDOjbwiL7wVKAcQVYZD/Y9X5j3gWXmT5dtBiEb1vMhJsXKB1Hq/P1qx47jQU
8FWG8uj5+lKgWkw868Y3mjVnLjkaM9AUf2JvvJpSrgiB3DHkyvAKJJ1Nn+zyQIKMnGcIyehHFHb/
rNXNQI45R3ZOMmjmoHPoUN8rlObAy/4HO4Y8AFSDkMgx0YuHBBS3nB5/Se4Ku2QbG9ZHksSnZ5BZ
JnaahleOfEwIpwuRbqD9BywSuKD9Rmcs1gamtaT3I39B5XB/BceA0otNB5JZGDL65D7OhGFyeKNL
+Vur3L3i8S6d7g4VKfd6aLbeVn3e39BXp62yk8H2dWwN6+iKpFdGck1BuHkZt8QvBAazhcFhbjd2
EpoB1V2+wnlQ/dR19kMk1N26nPzha89/JT7/6tBlSMfTFr+DUZDGGR9doQGEAlk25PW5flYQXM1B
uPTumtO6kMswYPJD9Yb/J3Do4+R6m4XALDTOPtdJZ4MCGl0vS5q0RiSOiytVpx50mNJM9/VcnRfR
0GzBPGa2Q78eG6WugA/NMX5ZVU+ks6HWEh0Axwu6ozACap8F36Anhf0/d034yH/VaDJwJUvRUSFg
tXTqdHdWrX5s59U7impB8tqBI4EI/cBe6jPGt04ZjMoU3GoFQhBFQDv+DIIgJHq/95V9q0EhGA/4
26kBI9Fk9G3f01nHVc0zll/9vBoLk2AzL6vZJXvRdvNQF9WaytCQFo+NZXUYFpJpSvjAITR6Ub3Z
9MukDOykW/bC2WV3IC2+j8lQJrAoNcyJiKEHpl5kUJtR3+cqG5r6zM9xuK5XGrASCICwJSRNIlfI
mn4IDZgfxT5YwK6g8jQHQwkgbuN6/jlENCev7EmFn9u8Pz9PlfbHFVOUFisXR9VZwDrgPYMCZuGy
YKlr4UJZW3bbKQeBZgJtKxUfu4LDhFhlssGRDE8Pw5QamwLrmJayY+u7iC13e1q+UT/SAhwXoO6a
bio3ldvm1Kqcna1QcG6WpJr7tzq+L0gP7GokAUg9Uyx84nzYP8/VPv+J7xBCirocwJDqCxBzbDXq
5XIPMf5oqm36p22ju72FFFJL9VXifsJw0ZdP1lZuTugKHJvdV4pBJB7hNXgg0splFhwtmw3pHnvk
/28cMis+6Ktf/bgGskQEFBnw2u/tX0lqDT4NAJw2UbrsuniUOy0m1d1XVtpEMpnUdcbzjz8RYzYg
DTuSsRZBhp3bhWBFUC9QxpJndAhPgqtrjo6/elr4gGVOD/rj38t45/rV54WIpmAjBGcakkyzs6Wa
Sq1fcRteFwEsZg1vXDBTL08vdfrrjpOuPgcDE9TP0WPaNX+xbh14aFT9ktNgO+Pbq9mIpMP/CIis
+QQ3a8bXJezXuSUgtcPw+oaO3NNXz/gSb8PaevBko2deyemz1F4xvHGsnWr8GQ/4/OcBhblha5Qx
UHV6Vrh73udwYK1flEoWvMwCUO2SwBCsUs+9xyWymv6OSvnK6BS0tM7Ox22CSqMZvOageaflNhFt
TGaNdtgJRjVHCPvGeCnIz71Ql22oTrcIvkJl3nlteD5eci5nmvjc7n5v7/H9MHJFX+N0MV7AxmJL
V/QAgNVL8hopZeeNxTAvOzhwlTPZnCcbppjZa/I94MHfniuxmn8UpTwve/QKRORM4BVEB/wUgiW0
LvnW5E0GKinvZD88iyy0NVc7WmSHlpleeYcM2ArA+qa0QRSN9wBtCzQNDBmoRa6nVe+9OsDEevEq
jOwX8w1Wd5nxR3eSdapXEuvUSmBgI6sJVrUbW4pURTq39h6XRo8a7en+2lNvqGt6N+HT1hOeQltK
aIO/jqK54/fa1wRzhlOLaXCYQ11qlax1Ysf83Q2TdEb9zQ39vAuaphHtvafqPOBmjeMBmpgxIqCi
ZxQk3gvd7VBf7fRCs17uayzC28wY70UkRkkOT8ZEexzNf5Vp/lHx3twdo/ZCtpL3m5CLXI2lUjnp
uRVUpIbSKJBA8/e5KfSKoscYccKwW6V9lZWrsx4RlixLOFO8pGC6bQ8VSiFwGW4/Ks/Y3dNLgs5r
sovgIu8E4HweIRydvFCrpPx6BbdGMHDh4bmVDW39i1Qu44WtOk5whhUaPo2Cv3U8enQOGjbtGfLY
Tu0yxtk9OuadNVDN2uUpAct+YvnQEQxxps1EB+Hzo4vuVeHsXu6UIeXLbufql5KzCcd+uNxlyJ9p
Lzopoi7a6B2+QiUeOUzr0qDCk7ilDnnjaXBaWgH+KPMWQ53GkeeDtnlS6ES28qXij0096sV4RRVT
tAWvtoNpSPfUnIjW+twe1W74mqRamC2Ph6gZKvvav3ZFJoAOjTxGmo2uUIlPRPr+xy6/rsFbKEor
wIj4DtoEr4qUumM5tggq9rFOVX0bNkMikrpLpBbGok6VcEDv9VFhQfdB7mpkedynTttKg6IDgEb+
7LChWXOwVeFGQk/wud4d2ZzgcJdQuJqOA2esEwHMqdOPiYSkI5y9ed02QIarU4H4fhEn9xg3QdXl
/vcDqhC0xNu8i/w8j90De9WiTxPZ5QExTcZqzByXLngKnUghvorYZk1cY90qTYbzpQ3h5hflSxoa
lS552GvQ1sPsVc+Od+Hi1cffNNRT0jwZbD6Xkc4+PByzXqZTn1oIzPEkDyIPbM77iMZpI44SQb1W
vFlpZFvTWeT89Zfbtc1IRq9W6GXEi6s86MbFKFeMEq8f/2dFenWSMj52trwN47um9iCpnBDDuLRI
Z1M0GNeLPFJDFLhlmeU3e7ozM70sdzsFvg34p0KEaQAmvedEEvviWCYeWSB2ZnJUT4NjYStMu9/6
JyUk9mtZUhe2JQyrjIf2HzJwuIoJwkfIBJx8bwljomg5u+BpB2OFNV3UAH9acf+1PBu5NkVJpDqk
wKM96UVQzyDIf11ABAMqmNmvRvdt32F46Ds68F42Iz79fM3vHJQ5Fjx61K8HIyfPWg1Br7qtH4VQ
QwDJ+pmLxKidpzWbcY6HQZ7SX0SjZxKAAH4J0l+i6mMhbJuzfJA0dRXqIZZ9jcA0xGNIZ/gFAP6X
iBlLowS9HNbVX4lr05B0W0JkTXrWnCYCW6ohZz5o849BeIApTXrlP54mmd4t5EsRXozaHTNZvAtN
yp5B53lOY2m/FwghhV1byMtAz2bEuMOLgXEEdgaHKilhTNt5NhjGE0jRjSmkJqogAT/2Kk+kDER5
JnU+ws2iMX+KKzHG53Zsm6ZOl4Hl+BfIETpfWW+hEXUa6F5BC2JRQvk64DKC7iOEzr6x7EkIOL4E
ERO5Thtd+bGlTm1FWyIFi7SRvoIYuNfOOj2f54XkVIWH3EUqALlFtd0s+SxLC74HvSN8aj4o2+U9
w+bntRqp+i3M+Ja/5uNsjFWldf2uetPfKXpbP0PB7aO/V0Hjm5UoOjYGdovLwDRsN8OSZKHqtwCX
4f2m6EFLf3FjcMDFjT3/DBSviEd8LgvtNBXtzxrPivcTVerSMKRBT8HhDnztO1FF/PHjdBOSN7gb
hOosWlK73i/K5sUMIKnBrILgCrBhbmlR2icj+xBXYrIXDmZ+tPRyetQCz7ihNlP+ux4UkNhkOJi9
W50ju4MR0xsj28Q1I8UFFcEDMrLbVm51VEksz+A7l+gb3DJ40xWjBawF/w+AZLGxcEBfZIsr4UQ4
p8zj20LfEZ0gjFN2tmsIJidO3qkUk0KhpO0RBR1iZgWuGDzbASpvGh8yJks8+xsiZ3vqOSNZCYpt
AFrpGI6WeFIWL30I3EFf705eE59pxf2/ZZglrLpY+jRv4vJA9Xmt93AFJ1joqvZEZeGvJp0iKKwb
0ErNgrKc8QY5ZK9EIYnOkR+OaIqOwLomboBCbkBJW20AtIo6VI6fKtSZigC1tRdLs4ymSgrYK7Ze
E+u9tGcs5hIs5ClD0S4uNej99/BrIoUStxj8v43Z3ahsLx/+py9UUTjeHSthdMWyFXzGgIeO8ut4
jUAbWYZEYkzmvj9nVcXKIumFH0tMtUXCf7s5AjlqDA+uJjFNJn4lDQUKlAcd6zUgorZioVMowPjF
pMoWduFvT0ZeFJaW/CwT6UGQECEnikoVuRqO7v0hvl6D2ldfbER/WUYK1PoYUQ/hpTzEtikcYDQz
yxI/CkxS9+DuyHIa36KYuTKy8R8kHsNnG7NwVM08rpX2RJBH2iL0grcLfuXZAe3ox0V0XcM4pM54
s6GMz7MmudwRAECsV1S2vopHuwkmoLtn5RUUOLfjRcu+Gyl4RWuD8PPiYD1hgwCv6QUfDvS735VY
DQAtX+dLG1hxw5V5C1VVj7NPe/rylcAfKKmQMRAr4QCl82gItYwqi07+tujNO/I0BFZ7T6uSXi1R
AlIUuuvG5ilbFeD9yWx2xFaw2DfAgQv0qVTMODtTyfVfynPYpe0HtPkt3XFFJZvWhAp0XXP0GGrB
3UOnDouGfhhsJUJDFqSpOXOFCJWwPtsIx85OE/HMdPW6n+y4bAlZDuTt66uRZUT084JliN438ZQE
k5plxAwUa3TC8f67Oyk3bpe3ySGAJqiUkpzGkSW9O66QyTwzlnVrQV80QpLf+nyTqxdjPTgvdLNA
DoCjpjK4h/x/VHqD81Mrv9FNxrCws5OIpTvR8JsizrGaegdVyTZne5bZCnBXUkLbU7VFubUJX/Sq
XkVPNUEldnugtDhxnqicDFzWGOySX6cueNWU3FzC6sMo3Yntb8oiRQMcjGgBtrz6zlJ/CRhORWQX
yvb2str1VyPPGbe7Zb+G47v7nz2kI9lSR4iPsI69xxVLOZm9S6yF1uPniAE+488jVbkzBRamnyz3
+3kXj+jcsM8MvfXYi8QMRsgHoo7ZEFB+Lzehd3E2X18NuEIi769EK/qR6yGwBdmJg9VLhLjICteR
7pbiZbG2KJDNeLlUK/GelTVinE0WI8NhxW9+3+EWGp0zfdvmNvGqiNqAT1HkaHkLjucpJtjd8tbk
g1k1YuYRf+RZmqbbRI8mK5NkiyoT6EE/Dl7ozYWnwH46Lo/75lh57ZzuQ28zzME8z6sOjN5R25t0
KTtqvHTwm5WIWHUTR4Q04ULsYa4w3H+aiKP+wY8n5MWcQOE7A7c6lXpvobMSHB23poi9nBOpwx7f
wLBhSZ3OBOHbdXUNxuoAn4PAWhOxhdHmCwT1IJxEB1Zk2q946tXaK1Gi5G7GyO9USFRb+C1UwpXS
08mGzbhBGVh9577QxmycZ4i/NWssjJ/+qDPxBrOKs98daSiKz5/5nwXrSmXGGiVTIwQXtDjUpxQL
2E86AdUpkNn9xDAuCzS4W1Se98//uC7XEDDwqh0zhF1VLgbdb1iUjMsA9Is4oWAg8yKDmSLeLN7g
I+JgNVz2GDarcY5aXSxzR1gTFXIv/85rxyyuibbHaL1N0evI6a+32pDkaQTg8kkf9UrVncOtbFpS
p6VA8FqyQqX0yDPaeKiDGx2yhdWQ+HAAZYEvjXOI96SfpHyEeEsJ5lnBb1qkPhtfe++ntlJSedA2
eVYVAxFF6d8NsKcw3HBJdili4l81bcwSA9uWKaJlg+FT2VclQsTWhNd6MjHgTm6jc9ILsOWxXxJw
YqJHHwOwhzTqq2Q6lix4xdbkakRqITs0BXvyKlYIHLv0tZ/MU2p/suYN7EYq4l3oYsHT+Khr4lhj
kUZDrTmFFRS0cSXrfmWB55tr5X3r0ZxU44bLJQe5oWji4x9teDHJ1/IThwpRJC0ogyX18q62SG+J
UCSgQote7uTlLF3r8hDqqn8W+bUgkGfZydYg8bWZAYx0fvCSr1U0DQSk9XdvScHEpgFg9ECr2v+l
6Ei769lQEMnOatLCGQUdW9k4wgYoSR2LZZnZZid9ByLyfHM5bttxDBYsFxcTM7yzPudChApWED3B
cz85R4EMzy6UcgAEXgCLMTtPCklsp4G9ri8PqXz6IFtVWKfykMQ/JNsopVo5+f9jORQZMeJ/0vdA
9tv5Vsv9FLsz584J/rgfkYV2l02pw9XltLHKK0t++QqBx+pUP5GaSpRtjNh9NF3o8vNXI/6NBZxy
C3hBFoZqrPp8EH035Dg6XA3ZvJfhLb4ZvK6GoRBfMCmxMtSLQ0jamlI8Q2oupT+2vzmtwAgSuDDP
rff6SenqCk3sKLz4pjWNnZEjF9MN7XFVPJ72KtnS/rmSWQXpYNI5XRnJMc1m98hhmmhSPtxFNoPW
byREtblG0JXw9IWXem1JvSUKi8NEfdbyx5j61YlJu97UrytIf2+HWzUD9MQl6U77phe6n9WLrxRX
n8LCtQMjMkpvxTr+US6KjrA7bK6raLKf1dHQ/HudabmZNs6tzV7c7x9mo5LrB0hrNl/cgr4F9Rn0
sfKAHDe9jS8oLy/WBKwopE3XeZMLuL+sq45O9xU2rEXc9SfM9zeHn/QDPt/wK0KIshYSZ7sYNt6o
Y3oCzArwM4BmWEKjfE8PAypgOuxidMoQIOzRD+v4msz94XMUPvi7KzoA6nbTYmDCK8VriBhg8yNa
+7hCQqWSA0pIMH7+kc2+Z907LkJBAx8Jz6XXTCWhMnOLbXvnmit1nd/9GWUEpnhuzbYQxGaTDdLX
ck52eMDF/4JA/FrrCLBkPH4UJP8t8MqUK1GR3B9BduvFUfgsKO661O/66HkhQRkFmdnyJvh+FE0v
/zLPjwFy0TANAktdlJp6gjKNFFWXemnci5IEm+dOzC/j9jb3pAkI6QSII9X5f71SOU6FfpGTIR1q
khV9QU6spxtTUA5JLTgvnlf8CNqEnGniPDK1/qKHcCIdeS/TnFjbRF9nBIzR8BxrHiYfphvWv5vi
2Jl++fgyfDBxpA5DL4xsy+FX+t2ccgMJIN1d0aj3Jaud8I//kCiRUyKEGbI7bn7ZqXQJBl/a9BeD
jLOFwSnDTqIQ1fg7nhOQ8jRs35Lz4aDHwQns/TRamd6DiaxPPOnfkfsZ5aLPDuKw176VxXmJ0ixn
gqXU0Q3s7X0jTeQhUHkr2QYrohSsi6BjiH0icV0HfF/H6E85PEbQbFaCHM+A9UnhZIOP9Lk+huNI
atNSnUbu2OkLU2LAq5icXwDE1UbCDpNU5VWqYs5NhndXIXQJ19KTK9CMBlrGf4+ZC5Pgq6t6iPuB
0vQm8CmnoEX2jtqYyotYkfrXhEtw4ycjXEp4aLRlZejAIxF0X1uURAFCwDMhY52lEN1ODs/T6uhs
d9P5NqB86ZkHQM4talbvQogyXf/NhC5QuUgkxnYzWr5ZqZZ9v8WmSZNJXCvMhnAmBDBucf2uiD4Z
+y9twKnbsQrhzZdV/Yt5Ub7MRnFFQv+pnvrf45GKDNPHeaMKckgf2aImhscu0b25o3b/nZM2PxCx
eKrDLk+MH/2ejarMgnNdig0Ubb4PuWnBQiRyUYBCQs4CyHvuW9PMfUiszuXHTD3SmlUckv6BrYq+
fD36g4twaSuzsAekD9HZFIest5WVk3fOl1Kwqzdo1WjQxy/TYUQ5ZlnW2TP1lJMEN1gZiEa8b8C+
50oMn+rxE6e5B/U3DbSSUCTF2OJg2C+UL12FVx9M4FUcZVnJmLSq/CeWT1+XRIrUwBuPRuih7jlb
nJIgLNiFj0xeFk4ivcdu63E4kwz5EU3KBEBDoMsLgNk5aPO7qpUHDCsim3fVXp3m5cW+15qf07FY
fMPLrvRBaWtooMCRg1FWQD2WEFP0efIcrHp719hpQGL1sXoN/6ySrAtEHznNhVEHCV8rUdUz3YI3
PPp/d0qo0XLd+W32iWbwQKTdYDv8VG0gcGl/1kJDDbkA4VGInjgYwJcAiuwr8OEqbPMocCj4X4CS
f3jWDczXwWGD5DsuH6RfLX56fOjjJvmmp/ZYggpb2NTjAzhiKuVzx8BFvLatR1E+vrZlZKhUjzBU
qlVtTs15sj20L8a1s5YzpLVLOhlk9vvqbecDMokpwAzBagupZ2nx/glVIB+NK0unbneYeXd2ZAvY
EepbMXBNks1aKMFtPpuUwjMR+SHOA5Q8tPww0O4ZzkscFxvYElDpSP5qkv5aSqhrw7wRUwJIH+8L
pDCkNMZ68AReI4hucuFECICU/OXicE6fvlAstpQSaYSf59tRh4tXFUVRFGJ5larcLbGFMIrviVI7
EkplKvZ28/D7xgWS0knsWoju5lHZXp4AmMRCV6tV+2NtY4dmcAt3p6PkyaPGweL7SBk+so9zPtsQ
+LWtA8ywmICBf7pSM5WjgXDrisaN3dG4vzcZj9giBCVzYWUyGytq6nGSajsmaLpHwzaFd8sGCed3
P55RIDDlaHLdjdtDTzLBBrDP3aBeUq/8CPUSADVXjhL38jNWfvwntIF4FikHtEMqFTFG91AbSV5V
Ip30IQViLq+udLcizwnfD/DXnyyIqYFiJEmnpGaNDvZMLYXWKkLw062fE40bBgTp3acGWyxLdB1V
of6viC+4Q90kVZmDFSbWKIPphm15s2WcYmruHl3xX7dX2ewETvgAMd9nKqaRVf+zty4WQOLVu6PO
4IYzIG6v+j+0vkphKTJkU3mp0H4g264j/AVs+PHqSH0i2MEQBjBqK0vrRlMWh/p+BN/f2evTsJ8/
ncYtSoJILaT8LnUVGkdz5HnBqFv8AsgLwwxvNTFGBaOxB+xWVAH91BmW2nYzb7l/Nr1lRwxgbzCQ
DbquiXD+J4isjvCN/n2dhi4IO3nZxqXi2X1E2eYkpvAS4SR2PPJkrkO990QmsAHYiqTVy5QjSl/s
wEghR5bbXLRKe51QEV9tsXp5EiVg65Raklh2LnXTxqb7MB5GRcOdMrAjaK9dUrlx2kIc3BR7v0H8
mg4/kde1sOhfzu8VvnvIihoipCry8RlN6rNj3ZuKviZ1aVni+xFqW8a4vhM7hW5M9NNf5d99bu8z
JrNNc5pAawRTWQBHB2kM30Q6UWVBFOihJYOOUUbUqYDZ1GrzfYZ03Jr5FtyAoi8FcIUrwO5ad9hz
03zhBTVEgQ8XSapE1fcW7Pkm2TIP3ZcjeQbPG972c44HnwWSHY3sl40CXcteOvCnxNnik8HO7TOL
C51PPc3RQFaUWjlg0Ph39dBB84ASXJ6yb0P6bE2cUVWQurwKYU65sejTQTbI5yGuP+/f4u+rTAz/
WHRZDL9iMWD6ilik+dhaD7u86Li2kwDErj18UKpeIgFd2wEdNlWCrD7ibrM3lxwigo+k7fd13auR
GrBvw4+7Q7FFrtxIhdUba/lWi9tNuyj+HNXw4s6VpzL7xJ4kFKqkyn2rItTOMTB3SZVMLi4enB6P
rPuAFqiqHIaynbymrgmoDZn+Gfvrp5NTflZB/vdc6W83AGYVvqkc95IBY+wkOsjC0YNo5dYEZ2BY
E+ci14tHezHNdm9b4nB5umBZOk7Ddk+gn3OAQWWsIl73v3cPVA6nKX0i16ZXDz934SmE24hgpOjf
JE4lCYNMK18kQzcs0d4C37nb5KmVJTiyTBAxP9oC2pI144SFn01X9VDxSwFHToSvuG4Do0cAKIsm
oFmAKUJiG+EoDE2Dmm0ofuoQJfSmhvlQpzA5H+h5YJd9esP52tSywui4YZqJiy73SooAV/CpOsqB
n3251lfC9JjDWrqeC8nXUZYsA44t30rIrucsJnHglY1esTY+OG5q0ybmtiXNcPfJ4ScqemhBSQ3j
8uAJpBwAFJwVnNC9NqgGvIiMR13/qNCgttRvx1OqG7pYVC3hX+5Eh19H7XElwbpN9S8yIZe3XmWX
vvS9+ECHGB/O/PvSizJ/EgsVvjCPpSSS2euf28QmeDUmhgiHk4b6bEyQyw8KCA+FpRzXmDmSNeQg
lC4NpeDyH8e+3UVUbF4q0ApVxB/w3I161i9Luy5RWF0Az8Unb1MZMqc1Gyt30lYvC06M56eMmW2L
BOGbzV/K5PBXtjC3WALDeR95aEVyWXq1pLRW+vNLiKpAj5uJEihNaOme7Z3GKgDDIFInZXaloAHM
RlqyWPW955U22Ax+Ggci9I/seq8p4mDiM5ZvS+TAteajmX0K511Zn2l+ABjOQp3QwhkZ1XM1oXFY
nPGwSrN4S7ZbO7P7z4NBccGz1YHs8ZXhhj1Rcg8NWj9pL8USh+HZD9v/bnumiJRe/uDYEJhocKEX
lk6MS+r84J9pfA/V5Th+SJuL7czNCw/FkiiGJa0pZqiq1tSwppY/wZdm+QrS/Uf+O6f70+CD1CJN
2QhVJIXIBgdcHDP7QW/rB2g8cUAHJJ7RpE94cCoNm9h+ieQdBRwyG891kLun+2oXBeYV+yA8IBvq
Qqnjv79o7UIuVbEGJjDD/oQKO3GpKyOZW/qcAmAR98KNEw5F70mpMLY0u7YArlY9F7drG450Eunp
5fwo7F3WY0Q5K0LkzZH5D5YIk0IbUR8CtwaS2BkqfKdkhkt7245whvf1PAq+KaKO2qTHOGsFAYP4
eKj4GPKZzArCMGA2xrrzRmL8eQzP8hwjHqx0AaQxrrwXpEX+SOLur81Ne+yXeqxFVwMeU7xwQHag
plPOHMLuaIEHJg7iB3jgRZ4tPl1z5rmuOfo0Z6MGlykdzvQbqRn26+KocFrXBOCI0SjfNHT59Zb2
XJg/j0IdMnf0FykeWcpIL674ncHkECOdfMI+uxiXJYvPeV5LLEyIrXr9AeOyZ1QTyEcgn/yn8djV
dnKpoYL5VPNCk8U/RfGtCPParSRNw8uOKzJbnX1h98BWCkhrOFFWYi3VPIkasrn33jr7Nu8z7zoY
CD1UcyIA4fqeg6fMf4wtLqmiDvV9dtP4VInExg/5iYh66Zb3tP072nVn2rrglEXXtkPx/s5nTc2j
tKx12v+Zxn+kPs8DM283TgYcD9VXXWmoc9XtjZD+hmZMDrzNCy15oxNvfvYK1NISIbdNAcRbLfhB
uWlO0XLUXc7TvZOgSFCLMQSqgiRHMGBZWU2CZmIamQGJbYyEidoYwMDDSehCuuRG2lG6Lp7NW76h
LUwRBo1wHi7dICNNnnYNDQTnlVFQnyMqeDsyMx1u1n0SBLrpGsR9n7Phk7JfCqQAmaz66wIWfLyl
SgpPhtEnxs49mtiu43BpAThtEv9TwTsLBvsNlorpQ43VJ0LeaJRwlNJQOEGrzd65TCMm6dNu8uny
7lU9SKwx1mvZ4MCjnCae5MrC6XYKQ9sij+lZWqKRs/SldnQEMkg16wqSnidmPoO3Qbh8YwraKqpu
NTvbUkLTRgbIduw66z6p98Q70iSreHd5nbQjZO+QXL/Sn2rqBiGVn3SmGQqQI0qK2qwgChAfPKEe
GdYE5/6wwxHfyeJFCWCWXxraLHPVu+1OeaAsmMEGa+Fen07jWq4dKSSP7OtiPWVdDRdCTgayCg7K
jTMH7hwT+8o96Mo2parCabNLqrQYFgebYA1/wtQZcnRHJgD97zQ3UWT2JxddbIE7whyezntNEUcP
eCWbPmNQPlcn04J+38dUMHF4YiZvaC+EA2YKaqDbvEo5jSSlzBm6AF0RDxCqWeR15zvvr22sz/Fu
G9EY6/GHEceKggfFKVLIEeP2T8OOfSB/1wDvaGO/D2RxMT7cuB7Y9l1Cbyc1QlO62DjZjwxmb2/3
Xe50nDRz97rMuI13mR3tPEqiR1ki56iF3FZmUREVhQR0c4bpIU/p67n3Oi5VN8FyC+MVr9Y4z24w
eT3uwfXmgjfVLanmSHHg421N+mq6bSo04W71fhk9ZDFWnaWm6rGg65VC80ZUd4as9m6YkoGR5NPU
nKV6rR1oxN45UX/HVfIeoLgF+ndOzM6aMuFv4soNUEMwnS+KD4SRuRUENJyPdEg1ToGX4cd/ehzK
VB3kzk8lWvnL2jJtMMErINslBhTvgwotXT5lReycCVs353aJ0X46fkrPL+DQ2NODReLMXYWXK8B2
i8x6seV8e/tKWr0leaQmG6Yz/+YDej2TaI+YjB9HWQsobbFxy6RPUnjaoONvh9xAfqSPSn+P/HO8
HZ+YshUVRFaI8J3v+1xnpJwKEOe34RyNOF63XLVuZBAhyBO4ZIoJJAs6HXcZT0t3gLbEw2147mvu
qBEQb/FoaqpmRTH+4OApx3rzvBKzqunakhvpbngCWNYKna2HD2oInPwr64k/9eBADaVcrT287WxZ
Cwymqwhd8ncaaXHhDZjQ0kFZaLIxRunyFK0Go9d5yQxUWX8MrNhxjZRgYFDACa24BH8NIrmBGq3j
tBPYK1A/N/H0WfBFkxtbxSX18/2HyM01JxeHslCn/cG/JE2sIj5ukERPqF9JCn1acC9WWY+io8JI
cf7v06EwT5k33+oku9eYgfg5qJGpAJCUjSoLniGISjmsFsUzg9ycQVqlkQt+lvK3zDFOJnN/nb0e
0hBRotrKfI6QlT4EuYE+26kBpVkRS1h0zj5jhvLW6g1+9xQLJSNw7XCbAI1Q8qL/HvYlKmnb8i/L
6DOK8J3zk+omwC9eXAef4uIRNNtR1GIxAiGGHgClUA51TLVthcB1+UuIjSK9RhbRSnllduHOo/Pf
vE+uoKo4l7NGf2iLpS5VvNFy14z5LbuJ7N67AIzsstEfyUauDRBx/aKydvURmsEDWz5+fpzQ990C
5ovsVmKmWjFH+EPragBV7c5nsEyasKbQ0HxrmtjSGHwBuiKwvS8cn9GO1qhuct2S/tcbg+Lbres7
uCSxmw9YS9NIy/7Rw4+KudA1hYxWJtCh59F3BJaQP/nVuvAYepgUaOrkWORW91uUk8EDeewfQORk
r2pB3D2m5U84V6AjHdIxmPUcKCLEMjaHyrrIkLZzvE0jg/G1f2jLrUsLP1nMY88qdNHLTpr0YGpC
dLXCgH4xPRtTboHgBilaELXdF9yBqh+4r1l1QrKkU49OplRUJDTcxxgz1AxnPAQLoBfrvt8NRR40
LzZQB6g11Taghmh8bz4wv+iT5WEVKFxIxtw7E9VKJ5otDevVReAxC8f3ihaYk8dRIbakDNY0bjk0
7JsjMf3H8HlTaQvKosV+4mkKJfNPHRSoghWXur72Tfu9jvmrNJROFZki9IqC2+F52h4l8ZNKA2Ko
3ZIvY9j3I9r1+AJ8xQUi9y+SgB7atI7xOiofyyP+KAEpL9yx4pyC1mLK6apIriABCXUq0NtqS1pZ
ck6obkJROmkQL4eaD9LwWPfgJJda7Tx05bR2uPo/XqsjOizcjGEbd3BQslFYN0JVPpUy5AQqQmo/
IHaw+mXNm0ufs+ppoATHV8p4yO4pnXkztCGxc0kla0FRquWl7ye3FfSgor94O7Qfdk7/WRsmrt7g
Fjxuy/5Bh4Q008CYwvbU1b2/oZBHgv6G10DAHCHswZu/YJq6Y+uHPoE5ecFfxWZiwh2RVWqrFTS+
+MZxnHANyFvF0FuGrmjTqBMpc3QHxEt2G15OzI4bfGcVjXxa9nJafWaoyDXTeJ/HNxVv5iTxxmIG
2pbiTngZVPvBTodnf7TrHS5X5NfZgbcc0gGIMxS1kWnqE9VZRynTyOopm63WKyhH2veLpp+/7tQi
ah/CcbwAJf5CozVlBaRmfgSc0Q5CQCgFamIehTGYgzZ4KV9BUjEUozi1sVGiT2hLOpfZCpOLGBfm
XKEAErDVNcANKNoLSXUmLlGRfb6byI66ClpP018nClXc6oKxPTDSFxC6gSWUs1Owub5L4mwWyBmH
1gQAV8jBKDMAi/49S/e8i6Z+VRVJ5o0VRYiBze0z4N9dj3t6oQ6ubgTSSXGUrR3ez1+ixycIR4+b
WJ/MSPQcaooue5ndD6Wqo7aRuWb5gTkEVNsf1i8Dwc5MJlJNClcAYMJVh2nYMT9Iuxb1InTTwcU9
aamSixLl5McXsXmizXdtC5d/KckJSKZ8uzeb7EQFby711if8GkYCFRfNMRYUJqBApqmcUIE5v44q
3z4hZS4BnZd6vaJ+CDeVSvcPSwKYeZHMtK2tNDQBwdwAXh5CKsUHDRRyyhxuyefB8gO/v2BsweuE
mmoAq8ArlXKiy7Peb0l4EUb4xHcmywsu3OKI6p1vmSLy5o8N1MM5521yXPqaaQ3VZ6Ts0bIFCHCy
2/SSmBpZbrQe5kBelSkIJq9gqLt4j+NRqa0S1n1yzGWWm0UsJBSXDLEoDC5f+U6X7iEWVTorJM5n
W7JyfonVaRsSst6SYFJT+CKPYYBw9eIfZR+dweEYk7GYwbktC1a12nDZM4BPK1Qv99BJfQLq+wZP
CE/XbgUSiQwDjJxJRVbnK+E6hUxW7egoU8AmcsPcG8AKNvUuTu+8ZTLbNceqcbZq73NLGED3h3QC
FGtvquVeIh2FHAFF9PMBdCZhJk6fSzRSPD9Uj6n+mlSw934FXfPdG5/Cb29K2Qz9zaYEC5fQ/kou
tZDQizcJcbx90YucFuOFdHJiDrzd/dDLX4AF6sf7r7mQuVsmQul8TO7aOFuVNIZk4715F09+RTCJ
2GF+nQY+BTUDK8whkycmcetio6EiIUL+j113dTbntjtPkmnJEY4cNHlPc5EkQVebjTNBNYbYlTi/
ehLLu8EcrHRYREf4WdozkThh798Xp5sbtGgyMnO/G12h/xQ1JKVL9hmOT3krUJ8QZEbqIOMJqZAj
lxkm8d+vWbAHdh5PsYRBUsQgb0lNKfEFE+b1oX/xnEltSE8fdUvheb4fdroPHeru0NDTCXbwDdNg
aypos/xYk27w98QL9rBuIixQmxjyG8q2SHa8squYXoOa1OlvCSKxqpcPtIxHh+5ZHLaGNqg88fD9
6U7AdcQf1cYY6UIx3TKmxFGERIXDeV/MaUTXIZVGwrHqCMyYKB11TiwiD250CyDll3wDuUmqgiJL
mA2SY6OHgjMwsbDlJXyBOO14Dc5u6GaXr4ewBrJUeh7iwS+IVCeNIUxp7qywKSrnd6WIaJLgkHQJ
pVKTnmrdJWgqbwi2QEUqwjYhCCkMcshpOBJ0LRHPXBU6qgkGgfVf5aklxfpJ5kWpHIjVBxjKFBOF
hmoZN8moAiJ+J6neiWlCJiz426xIcBB/IPGzEGfbRkLsDnCkfRBK+ifl/bKhgi2fCuqG5hPGedaG
jHg3HEa5qrGexQ2xipMthKhjqR7gwO3b5MysajLTgSx+tsWKdpWsAI7iAjs3h3po3LvRvKYIGw3x
pSukTbwd1ZPSnI0IWmoVGxw88LmW5k+a9AH642KnSWFtkFbgH9ycZiv2IXHYG9p3kTiKeyGxOIS5
Fbyk54iEBp30SWJCZxikWxWXDkE15S/bKdkGhX/3f9h2cLecxjkDk4lz9UQCoDhhzhJzfrSqFcbG
IybP1+v8lsqpatf4wL7HzvyG9uICDcQIo9erSP9W4Tmf8oaC3FBPhP0B8Lgb79I8qKRRDdfrAzxQ
6KWfB2H075AX3FvSiPfTeDIlrF+s9vuh3jrjTyci7TVdoOwqZOmKHDoYs68ULQXw3ABQRKOPWKQH
eERp2C2vlq3q6GrK5AEv7hJj9AlL0G2IdwM0g6RR1t7+/PhMvzwwFlKyhD9f1kmT/MBklYilLOAE
O+jGqc6pXvuoaqM0upAe4zDhTtZ6dZWS7umk+kl66lMZ0Hm32oRwwjJYVE5fFTDHBltD/GtMzYu+
MVv59qCXU+qI0100UrBlZ03uxC8fJ1nKQHuETNlWlKqcgf4ESCqm5gLlVJdy7AT3HZ5JHDCzotLI
FlbST7B7Ye42vXV43DYM63YHM9PsTsRe7G28ZySlZHzxhi0NhTe69oH6iuECPaa4A0WkKoiK6Wcb
L2752maChrwKUxyEbENvABud1Xa/9+muI1UKRgEv/YsSBlPuBrawRHvXgh+jRgGesC/jD1nWtdRN
NE6e1itVMq5B21ge/9B+Fha0BQ0mxWJKiZ4Erp2Z6gYFBTVda6WmlMlg8sfFueGBFi+j+lVOPcAG
hbeCzrXTCi0kSfdpxjoZUNE/P4jcky9kBJC5fjVeBYWshh0nJNu5vZEJYAgfO/B68n1Gs1622a9/
BN9yQPPBnM3vZZZ1PwMm+xZOkZPmr9FReaTggpKF7Hs0feQ2UVFDFCZeRLCKDMYa0mqvwb1fBVbB
1IgedeMkLPaaclfkCLZsWRuMb1aLLr4x648P7YMJW6NwGVSKa+VltsZgATWE395+GRwKtkUSPdGu
VLLVED4U1kNLC3cLaDIeAo8dNgcpDviVAm/ZFKSaMkFYGcZvD8SljAqnr/1WXAcCEwNxsXx+y0JU
6B9WKSM7ftDyPBhSQNSLmVxVpXpmT69tYDRX5mxf1abMVPXZ6fDoUuvuGxLwUcev7JgL7y1iYw37
D4PHkaZw9K2/cZ7vm1WCiw0fZXe28Q5ZDomhGg6jfSaVOZvz9teYv+T8PvAouxfMTc6nU+Jz9cO/
S/TMinxyxHgSbdLKFDUOytbJXx7uXYODl52PgumjTLPFzyvh2JCwu1Bwtz8t8p0f8IA4bRRqUUwq
emRpVcjde8jKw2qMpQaPI2Yock1yADAjaBbgtnsLGOEzKfBwAGw4mD3IQFEoQLQHY2n6rusleUrZ
dR1ZFySlx2y2dyaSiNFqjYiSe7cOLf8DGOBvRr2YtuUDgT7twqJ+y86IaKKdnIlyBBiMcAMTO+2R
2xmx75P86zmqQP//IuGphnqoifNwX+e6rLtvfKv/XEprxSaIrtv09XFP1l6XHGeAaldhf2oBnsBg
s3fc6851SWT5B/rKdXoGkA7+W+jqOPbfa846A6m7kmwb/yg11Zhl1rsdFd5Y7uO77DgxW+EjZszg
jNMJd1Z7P3Ck+SJcLu2nb5WhOgVRwCXN2xa3tYZlg0+pxQZeKuWI1F5CB2tWk3Ob0XHGdR4JUbiO
dJ6k/ptiopOKDmwsVRTutYjIImLBXAoYuMDvQf+rcJ155/oiRhAu+zm6pXFOxjnCWb9Ax7Go4Lsr
ki9yU4JOrvhZeVn5+Hh9oHNfdFSS0EsQfpEGCZMK2a2VzVzEOCe6ggxhcdr1s4zcRgpL9s/zqTQm
1fNXU2tggJ6oel9UoBCLjN5OOdOPDRfehNHQLFkFogEVQwlaexr659GG/vHqj5/Kj8P3uAhmI4c/
9YR+X6AEeHiD32k/GItmZexE9pkup/yDWr7627Ur34wQ/2ctu8rzoY6IOGaaszTf5YS2o2sOVM0U
hbtCoSnXF84PU4Figf/vw6aT1P+nfibhIzrNv/ChyWjI0sAuCGs05bQb4ln6T3+AVy8H9Y8mOa2y
gU7YQqDQrCT0qiVKL76IxIfXgOXiA5+Z+Tz32jw1l1zTFcOW92obJtb8ZHhLs1JxANYLcI2mfXbh
z91vcJ0emCG+j7bUsCwpnd6hIFBglFbNvQd7kp9jSwQ7z1ayZZBlihGO3jPMntosG3Baag0lb7GS
X1S35np7lmGbQ9/X0V+xiZcm2ARw+av3dfq+fwQi8Zk20TrBqE7N9NEpgPBSb/NHNr7MMGRdVQNi
ccGAkqmHECpOPeq1Hd4r3gjgffyzRwKJG3Qt0xm5oKFsHcq5mdOxMnKhML1wP73QT/CMYoscpmPE
0+pb+VsGdsjWbXOCZ4FTQ18ry1kBQmrn7jmqDDma3G46258cFI29pX32TqQSwDQteMHRL4/XxZ5N
hIHia4XQVWfAI87MaYznCN/kVNTC753RqnkOZgXb4SiIvzcxTRIpEDyV4FtGac02ykaUAFNGqZVS
XnqN0KLlfLX2fHv4dr2DI1c8i4liiKIcQ5sTX0eFJnvKjK18onhTBnSUWOu5dDSeBGTBVp/CpdsG
8L+lGQ32ovKIitTf3sh8hHvzaz4IsBbyNQmk/hVnxHJqUL/+ImznKnW4M3WiVyi1V3mBs5iONtxs
m439LxXwBdpAKYPkYRBv9dyc/abKJxEPWtW56YF3jlzBcpaYBM4zSHbgqTWE+Uv+4POK4NkNhWsK
jl+yloCnqkIm21cTYS8xZg1Zr+zRiFaLAISxMhaClfofBAAYqFPkz6QaHs95S7l5opqoD3ouXKQe
CplwPJN0zZvEdCLR2yKZQq5l4VKKopOyrIwI4keFyhgYc3nhDwsHn8Jvm0yRuc2woULdSlwxX8hh
fWQ5KmM2c/pnF+roSIlTXtnylYzZmnfS1Fnu6ylx3aJoECv/5bnzMEi4nsKYjbptH1GkZ6fD9Mc4
DFBC9Nft/d8+fVOpp53skFDr9c1qZVYVn+A9qUDUF9YEzCaBBDrAYZL14ytMHOlT5EAYQKs3PMAN
Vp6TiOYCDWFjoEKWkMsPuRLa9Roun0l/Eb21ty1mVrnogi0Gkue4ANqqjC4XbSnZC2x27WFDNbGK
R1CJJbU4+97OJp31ljzVG/DWinKnIWXiJxZ2vCrbBuZXMS5drzcu3cL0dZa1JcsPKmEzOVKATemV
Y4kiQYgrG1v1S0qxjJEBhzQQJ5rQvRaFjSz57gmuYfH3cdQaUolNql1F+dvfigS929Ma73H2EnnX
avz1j6fYvXTt0vQW18fFsDEqgXfCkXEvhftCgDZE13su8kI9kCtG3cmKXyDCMX6T4s3dFyOCh7Wb
E1N1/ygeTWajuFV3TdmdWxcadJykoyBFZAJHUIZJVubVxwwilLVJKgI/XZsiOz6JrXu2ABxpp49z
LnyW4qDJltD1MFjp2CbpuMJL98ibbqJJcgh5PTREI8kTDWdOZmAymK1RTYWbG7vQd2f/2llRteTh
IJyQhLIEIxoYIxK0lpRlFbAQpkmmkd/6mNeJEjK0Tut4XBbwd+pcZH7zJpve3PEU7/OnT7XFJbbb
U46nxYsijH5GrqYIibDvM87RGHztAzOQ7/qvn9F0YvLnkfjhB7vwN5fTmghIPjf2Kjeplpps4hbE
sXZNOJZpZ7WI5e70+vHxSsT1bi1gMGgadNv42LVsZRNi/vghwux9TpBTtMgLZ31QaSXuqj3uw7EK
VuljNd7FVBAwEwXKJif0aJHOX0In2rUjjbZEF/aHuDOIUxf4zBR2esgBON40Mb+QThHfSyQiuMZZ
lXcAFgsPZDn3o85iJnD/oDtzh68UTgtx93U/snpqZAgFvAn/pEkji8LosaGgXXS21WOq3s67oeQA
HVOXJt5P5AF8Y9vQfq3aBrqCBaQAvBAcYxt4TDv7GU98t9yJ7X8dpCEwZ54lxduiWcrpZyxDktx0
cuAK6GtVMp8HiLSUl/hJKX4DYhxLeUYcFGFR1fVmFcyGMoNVdXuROBMLlyqZ9GlNnM+nEnfdgBUr
emicxNWTh16eZ2l8/dA18FiOvWfS3Ldq4BeCCgtiaWwW/A/eUJZ/GqeE0Gh7yc3pbgYwLnY7dp1G
g+6XAIMYzHRikiGqkKdf3lQGiTs2TQepBxWRwJbzBrPBPv+VotfJpxBBsBWalcbmPRBgKQ6gIeQF
mZZLsCNBcfaf9WDb+T0NA/Xruy03gIWvxCD1Hqts3UQ+9/bRNLUxis9jBkbcUvGeIzqS+sM1poBm
qc/siIrhC8JNbc6TPT2iaKabI25aA/F9ESq2zklnyh8zXeOWKRQJXK/Rbc4FX5mNaeaudSSSU6j8
v4Lq1cdsK8tkE5L3ci3jPEF2Z/cDRz5vA5GKBqxjaZLjEyX12kgOnDkR4RDmhCGzVRmZK2PseS+L
htfnzmMq+G/sqXmbEJFGepDTUSfYMXQVu6yf3fa8IlDqeNQatIJdB1+gMxR7jjk8GJ6+g9/5jmNj
/nbsLdazJpj/lYJunw/7pOiBcO+JsjXX29JJUNMaPDKopfS7m/SA0/tq3M3v2tJYs6qCHaVLw8nB
7p969CBa2Hb6atrs92kk2F3MYk6wHaLixDuUW+Hb7CnRp8Q6f9+BrgINc+St46HQ3JQCFPam+CTT
1tnjOkbgkryKb2ajawkjoz3aQKHutNEZKjmUkDAM5L1HLpVnRtGp05UbmB9NMeOU76bfNqhyd5Ve
1RleM2Ucqj2GrAhCCKqISJAYdDT1+MrP0ZP9CsgnkklX23Wuu47f4d0+vL+XZGF5yaUq4l5SGIk5
Ur4Z+hFoWTPfi9y10Dra0iuzG0LkTtjam3zRwLWxGOvC0cTv+F2oWO/MxPynDsokJI99WcoPrylH
0TpGm9TVlMIv+fnbZWS/R8qtHi5aUD6Rrp5NEJo8TfLZa3rx3K4aaQ/63hPUnCqSXe1CB77nVmrb
uuXWdAV85MzFQH/9CuBM8REc7dSQ/vx4xXtksHGPn8SbyuwSNcvCZ4xug3KTrIaN+CmhMQ4l/Fo+
9JqcbN2Eo25qKrjRs6jNXamXPvgEpaz1vhlyqXD0wdt9g3mF0B7XKTEKYWCh8fQAoigSzEr3rD7Y
lhyDxIP9yBaN+mLdU4LwJsYnFsB8CekrVBcNLcVpC0I8fkcBWOKR0MbkVueyjPqc9dlr+Do1LJyq
Gxpab1Po6LpPVEejGm2KjRwlrj9twYwnMfw584BJTuYXiJkb0LUMntVvT0tN05NPtYSgm8xDIo/3
ft6vV7lhUyvyaAIbO4SQD7zfqQCcD3HnsazwRhaoKCJgvhgAT6d3ywP7OC1C3AbJ8lJeeu0ehmk6
vUQMGgnJaQEvFpufAIW3pq3vsDZpRvwYMDXkECbo5wtwdIjwFBFxyuQB3IVYmD4oR4+ta3Sx/1GD
qtqPzzU8MhlBpqtTe1dqB9qE2gb1gAfAdZWVdD7WA4HM+ZtbCaFUs6Uos8QQBWeC6P1AzBHED6pS
YtUYMRhFFwzaavVxQq/gFQ0sff2HDOKtMQmsz7OJzhUwLJjcBxrsnVIm3f8xPqpYVXCbsxGI5iul
mJWkklIHVZ0jWrCzS+OoshQ/So6NSsVuxeTvNpf/0U+lvRXzLOghqdZmMnP2h7JOVmuOTWykg93C
P3cxhjHo9f8xCoqLaPYbQM740Buh+jzjwlHDTaFBU6eevVlKi73xUhstShXagkQfayhDDuGqkbXC
xapLJyPkbefXs/RDhAqkZvMxGylC764onuqHkxLTXHLI08v0Lv/2APKdPjl9QgPx/bQKKw/7pT42
lJkx7zBaucvNCISw55zjMACATABf/i+iOcHQPDHLTX07MVXoIcpjREN5oLS+JlohJdSkRLApXIrl
Oke5lT28YmZCO6OBqYC+yVPSxarFja5qGQqDkQOuBe5zxqFz81BuDqmRMKubPqy3gEw5AJ4tyr8h
SyJG91BLuDrkLLF6mKNno4p+/Sijh5HiKgbDcXU2TvheaZsDxuTOEHsKGLvEYfWo5ETnIC+t7qqH
ZN99apkcyg6/aNUhN3mjw+fNYGheO+4taSIqh4vv7xi8t0tijRmHudRqvdrvxsT74hhjrVC/ItgU
GbuFhO61Lh6z7FWPP64hXRnSSxmnAVPMlCZhvxTHcdamPeJ+d6zQI65/SMw/o3MOGDhChzJ8cTRG
7Cvbv12Uytpzn/Rv4ejgVAhYyy1bC8RGkKHybFsV3D7YlvA+8DvjM1x1xSi5hp84+Kq60/s2fN+q
NuSrkBRkKApdr7XUKYWuc6JCQZfkdafxdhlH8mcDKktCNEqf+zlG7UwTv3wSVpniIoMJKnqiPZS/
dHWPCqXkRiAsyJxw6SW4BtggPH6j6tdKQLkJQPEklQKI7M/RQHireNHmKrQvSw3a3s2PYWxq4xBi
b72ua6moE/cBScOerPgZ3yLAzlJaFl9I70stJGTbw8Cn5yPnqPnmAsMxtGDBVPE4AAgF9A3XzETa
8keqyejcc7xm72C5rz3GBmFKtKduWXMie7+WqMgRYj4rA6MpgBqD8JLrcaoV9IcvsPIstSKYiUER
QX0jFcEs8pPmAptRYajeLV8rFAgDUe38k6aslkI9Rze+2Jyfj8MVTGYcp3M3/hMBHCcCvmpzSMsP
6QEV6cOXIe8WFlVgI1DIlnkutEGNLypTjLV6tnc9HRSuKIugEuerZbNmpNsfRL2S5QV99kwKF3CX
qUDBFLT6gNHqtuHAnR9IpNKG4GjeBcgK5nLj4spWj67WICle4pVqXtjPaDcqnqqmRC7IuBLlML9j
mU6OV0ORckOvBUrI8dZ+1zrLfWPdAtYvmO1wlJoK7bUk7x7H0ZywJjLGXgUVPW1w3GehvJdWlnCS
617EKcz1eZ2rnSliNfDEjgwaAUhv6FThAOKLrQCfrZ1vanjRLCf8I5nIuZIVFpSXtPwF1XujewZp
n/o0wnF3ZPETwDq376UClB39mFuVSgaq9lcyLc1xle8l6PJouWBtZ1nucAWbKIGTkjL6Uv/KlnoF
RgOV3+qI4g1/RS0XLLMzZEp4uGKbWbxiIpzIP5m3ghjIDZgoI1q8Naez31Y8w1QnuFw3Zl1qn0WN
eQWOw5dwDReMHpIruRH7J9lxsAJ0DcSug2lZpNRh/TiJOvhjOrUxnGmKGa4rrEbXffZzTaBo8wtU
02rVa9NR6lCpUYAQSXYOjVZ8D/f0Y0TEKP/ixp2D4oGmopvwxOWVt7ipy924nErOthNCOCqDVFLK
OlJ/Y4QlQbusP5/aPBB8YhXKiELhgpTxE9pHnq15K9IMTNSecJmTNhg6bl9WdoTc5b5mVS1TjR6q
hzIJK4sVziDJZGoXpczDnQXLeskkJG0un+9/XenX6svT1wgZiCE6Rrt7lcl4uW7uy/SMwIHdq7jI
LdAcljSBy3JR2XQW7Dii3l3/5pzh30EVwVqqySqMCXW/NJNWOUJfftMlPDowxNl5qDWffrP5Lyuh
i3imPDrt8Jk5cElL2565dTGy5b1Mv4weHfnofYSzZbJs9uTOXttEHjPgZ4pQzG48EqXhdwyBnfU7
CntixyAXBdoC6g9f7fZsyV2QMHR6dPUXcqpigGu9B9E6+KH4JY8+/+PPsAXeDSx+eHk8PYjGVG72
zfbfElcX53nTmGCHQPpZWwGB/NXKXRA+qmv0zOLo5JRCEIunXXPcuM5UJzqLoBSSFheqqZDFYMww
Lz2Z3DwBnA/CGPdcNqNs3y+HZnjaR0xud54s5CJ/iLGcgaHekZcMrXA2+ce2J7bqE5cMdpTR6IUO
UM2CUNDWYxJo6bsH/lH9hF8B62R1ANm7fFjOPZe8VqlAKVm6d1FbSt15hojgtellu2zisAmBfib8
lEq023P1AtjxpbVKZ26bcNnbo9oFCDr01W+qDMi1Fmr49AtLjUXTJ2rxlGWVQ/KzUejok17l+VKe
FrJ+3cnj5ZrIcMvYrnTNFexPJmgNfi8PBbajZezJj5VTXGFWU7wVbdq3m+8SwSG7iZxBW6COjoAI
JQ0iCLoDEzKaDaPkwtkVXuU5DO2LqX7HeUy+P4WReVfSau57zuBxR0TGCNQq8sDWtQxURLo2zr93
bbkiE20mdfVsa+f6uWo4G1qKH7DZzi2r5ICFWC5yQCPgYtM73GDv8t0BiFIdbZrzFgCtf6wWUWXm
2vpIFSd7Y7xP5FZbIp3q7JwpBB6McwUqBF2N/pt3MaFdqKbFP2nkD0zZLd20Ra96kHd767O3jJwC
Y0rBMTS0krkNBYMypTyRbo2/lzdCiBJTfkVi6DxiPXmSKd9jTxpSEZpOXDcgpfvNX52RlUqr00TI
psx17FokczBCivUagdet2jItC2MC9xLT7LHi0g2k6x1JlQL3dQX/ilrMqA/GAxoQ0aON0ALpK9bO
Ks7LYJ0AeZZGtEZEdrP+Z74iBSZ8UVR19wBlpUBEUMSBW4MnNFZEC8wB8l4fB7S2fhjo5GOxH1OR
AedBxyihNsIecqbKG2M4ULD1L+zTYmBRIS47DIHWi3lUbMma9oDeqawTqMa9yMcQvy+jtBnArCGR
QNfNDeBGX3GZYdOz9Vz/p/zoG4iCEpnxw8KUbalryGDbEDHQTdqJbgnprkZ1Ut8uGZ7JzIHjMVv4
O2oBLSD9OevK3ry3iC6qhDAzLjNMC6IfjKjFwNzu0ZWc+UQF/ZIRjTs8WMbbnN5YGOx3QO28890Q
KyiWyCuX8rehK4Y+LBt3JteH+T1l9TzVeF2fu7op8oqnjvcv+tEnmISiR3zJyalbsjxiwsheu1vb
qLP4wl0TzQqmlVzJ+mGQ+O/ZualcQl3EIbEEjlth39jsEfNmmbYAjYsWR0tU+P82AJAnRSB2pcAB
WH4AvmTgkq6xt52daoGTu6tG0zUdCnfjWNLPGMVOMHfWT/K4VyrlHb1+T1ex5dH/47GNPEN+bwqg
2p2z5mVWL+e1trqAwaXnlgZ/DGvpHn1+lQZFj7PMsfi5i2DW6mJvzkrDScatklPK88C28KUAb5fk
Y4B9K4TMzS2Tigf5I7vZ4Kv/E5zxuStMvQLyys5Vq753r4n65FmFu/02d6k+9vgP/cVlmVuzvmEK
pbcfzBaYV4iO9u/hkWseYtk+cZwIl8FEeTsjmfgNgnSTJ8+707OoTZ4dU4UqgUxunECgZ8EL0/Sw
az6dHqlEQGv97QUXmKl3UE1E8xSHZydSuzYRO6+djPntG4ABrkIK52L6Jcl8ItjRY4VNoZMNMrcF
FLQeNxnALKEFzb/ZO61XRi8f2iHjxYESBNW3+icoRKS9ja5tT5ugTWkpByKqf/Y5sf9k+0zQSav8
wp8dec2DW2pP/2lqZlY44s2vqTrRHxgtJNeZF8d/kC1b9m1Zc/fuUxO+ePNAcB5Z+FCxyFKou0Ga
uDLWzPQbNPLn45Pfil6Q61mF7cwg1wpaZhjd6htrBB+JLEKAKIx26QoB6yGvn5/j9nXNNxDn82pk
fG147RcprlkIT27F0pH+XW8ZCABQuiPfvUl1zoe6sCQRLWyppQ5qVYH6hdtDSxriYFgzvh3EVs+g
TN+Ijohk1T7lEF/rhS0ntZzz/tCyp9PfCNKb2dzapKk46Dtx8wSRzmtK14NXxPb9gUP5ipoG2m1Q
rkqCbastu6xeu/nXrYSuowf7yCVRTRNyT+SlK+M/8J7c68BENktdRvLdpWTNqYphyxY2byNtTfLz
IcaaQJuw6KG31xOcDhMkk4oE8rOoUHGhw74ts3OWnWcA6qDz+H0HHNuhdoja0bMjOajJ3yNe0dvy
LiG0aVyY71Lf3xymAku5JLSuWq2JEY5v2Jx+FBF193u2xgxF6Fvq2T2UmdMUG4L0s6Jpcf7iwnWq
Weg2c6pNJ6GkjioAogjY+CvTFJiJhO05NFe8ENptcsT3S9bP/0I1aMYTf3m9fzvuxYkRD1d6CyI7
z2W4e3zLrbIBICmKW6QTRCur3hJwEqbZpQwGTG/6xzsQqDjlBM9f0bpZXQGD9KedRJ5Hd4VVslrh
ioQlOCzpmrtPbLM5eBQfsk7YnzzfuTmgvkrCocM2tLSvhOn4aUqdQYpvI/pm3C58RlH9a544cNfj
iujqU8ZtfKISyOoJqGgjbFJnLbBqyNEJ3REuLViVPSKd6FBkGuefsv7l+3yZEjJp1eruxtSa+bCD
KdMcx9IDAABYc3ld4ZIcepftfYCNP0k5wJrCgs91yTZIvAYSfgNxbPbUl8MygN9O6p2JeeimZUz5
41b1biQmgv7DA0OVdDbko5AosWpHNsis1ns8JYHJG/3E9o05oTkSjwIf4nMlw277GSz9JChPQqTI
i4/6kUzGsKm3y6GDZ/7Yl3pdyUEtxoBGouDEbsZiL/Qiy7mDOPJolc1c8FjYbKmQkzm5adKM5SRR
+F+WKmaxHBXqPFE3aqdBliiacDogiSY6CbnZFYzg7Mtvb5fXmGVbf7OitxOx+ywx+56HBzoUVEvk
39PTueJLLEsii/WhgdLKOJ+c2IiBub63bGf2Tkjo5KrpxTLVnW4ja7awCNUeDSlceg0Fx3xR/5AK
4qA+iUYo8R+jIQ6E6Uy7Y1lLoy53n3MH2360z4hlinkxnulaDlXQWqRNExpc18IyDQjPgttPzciW
vmFqK/Vvy4brcUPjZ6cPMikTjljCV8vsXiw6GEwaAn9WE2smy+Nv6v/KCyYHXLDFPbkF6PyL9PTu
xTMalnfa/3q/S4f4zgqM5KVq77UMXhuvckqJ6Qky9atgb47VJUWn0XIuhKI/7itq2vAkyupL36aC
ATE92KIc14PavelAM3I+kiV5U+26EWTCJ5sJBIhh2HUojbjwW2nAXDyMOHEG9WQYgNyKpD5sjCTz
QG2Y72lDY0blSRzqc9G1oofU7CRqiyLtOQFevUptdCI/8BguzB5WnqHcYF9+qxWYWRbS4CqlPY55
G610yMuB71tYRxhJCSHmLuOZ6SSpUDFXLjJAj9bKmxRCpcqg1dJ29/qoZQGZ3QTUsX63EeI4axkZ
Qe4sTOmtwjoUogxlDquSY9BToZZGD/6rBI0Jtf9UIY3kwxJd4pe3LjABcHphVMDqH+JFPZMJDw3h
9N/xGRAs2BL8tvkONfUwA75VSvLTidui5rXCsD2UbU4gkzvKwplwkV5EOB1YpPeLMZTaMEvVBCfr
E94u3op1oY/Iq4Qk4eQNePXaEfXbCRFB0MU+krt64tXnQtOry0lKFhRjdjevnsI80qW6p9rWdl+Q
53P/5LCOm2OlnbdLDu1RV03xfj1SnubcFG3LMeS8ZQu7J3Z5cQdbXVYZ+uSypct9pQSC+ghdZbfE
bHlhpnpFmF0ZeiHl8ml/x49xXPgh1DwzuDMIlfRg5r/hnlugnPn8r1H+eSQo+F0mMxsQTp2CYAF4
L3juupRoyFlNNN0utNudLnYDxCE4bZPbayGQwogA60dgexrPmec2290keJqHDa+vvThb3SAy6z9i
JibYTcGwmt0LQ7mMF33ux/IkF5nXdBW0TrCixjp//WT/mPQXCrl/wm8ryKK7ukBBl2EeGmbe+MLn
mUkJ0Bak7ExZmh7+9qTwoo8SYWdkNU4wseS7a4vR4UMU+0OWRKCip6Pp8hIHyVLM4H4EU6GiSQZC
QeEHGA6Hkj+Ik0XA7B3FHN+m23rVADJsP8mUY3UpwNZgSt+oFpak/IX0/rSPV7LdTq1gWEVWbUCW
susCFfk7auUfwGukwOs3QGUiN00D4vKHNnQzT9bMDyXgbc2RZ+Jq7Jo8fcDcO01/ItAnW2BmKXHc
pjgmPZ3YZWvW9MY/pxyfD4F3sbNT2TwYJ8b0LfQlKoU/07Mp3K2i3CID6MrwbG8Vuv7eMELJW57A
0SJn1qSHQjQyjL2g6rGE7yJOgPKHCDVRsnjJJgqCVbTrhq9OTMhHnbTr6SdORPZMSIhpIRXaI4Qi
HC9sG6arRF4IrnrOkIj0/qysfzAhRzt6ou4QJdDXLEmNiPlpt7f9ee/8g9eKOiGxUZUckkvfRwy/
8vWnPCY+OJ248WkusZ8CC2ymo8Pao2XyWEzh2UJBtvV036SYhWd3ov61yj3w+FQGbXjZN6QmxSlN
1iz8Wdv2j3OPhwTC+3cOicByt00QzMRqejup8SwIr7Smb6Zb49o64n1i5Bqi9603CNxO8MwjmF4i
xfX8x4HkeF8en4jAtnTYoQLoMGv1eplGIE9iD/JuQzIPI32hZC1G6kB5jJT4OoCyd8HkF83K1z0c
0Q96CQyLMF5mU74427iS9T+1E9/8jl+SB1o+Al7iW6sLUBUlUclFqwahB91N8UOZajuKItr7Ko4a
i+1jLCihCCHzGNptXuU0qIDUX09GCQLbz7Cn+zoB/xJ4LL5bTbyqJlmM7prI+T7mWTTvIWc24kEU
DrqkutluwDgE/fu70j6xszik6YM4Kq/LEU2Ojyk1Gpe950TJki4IoL1OxuDihBI44LPG1LNHNPI8
euhgPQzoyX2LKXYnCRgoaXDZB+cgTC1yzcKUUFDuen2LHXCw9hCcZXHPXP4L0yPST7Z3kVGZ+3gt
8z3CWF428UgQ1DToHEox004CXhKheogGgc/YCLFuHELL07pasCg5I86Bz1vhXvmvuK6rGp9XQ+wk
u775AmYULzok2EVG34KnFGacJOhnLH/C6IymTIkMnNBBcIkZsigaUCa61kYa8BE7uAAToi2/bxaP
gkbca27aZde3lvE4YDIjOLjqnBGL50dSznEp6bGGnLR2XUhkViQT8avD25GvvmPteu+3+cKQjBp4
ew0OfEU4JPt/fpLzT22lbj+cLqhXDhiEQfmjyM/xrAHnLhZ0tfgLqNk0nnVNZI30Y89isiOr+Yno
ZPQMV82qntshU9iDZzDHo3P4SVdyotZBi5eMyrRtqRqXYfff39I2tozfpMq+R+DQfukysvRO9e5S
aHEkhkszZK4CR5nwbeMRD8y/E2VCY4+WsDLVgLClENZC1XowTsEERUfzdrZJCb+pEAlmIciAOeWN
ulXgA+sTPTsT7LIgmhL2KTIAdzz5um9Keo+kyl6IwbiJOs59MKTsEJOALGawmiKnAYly06ju/KiS
QbnEzBNoROV7HcqxZYGaUThdZ3XQl6Yyra2eSuqgPXlXVaetCufwyDUZ31D2KIBL+OII5BRloyr7
5FxVVkb3sbW2mQHnjcny1mMVLuEqhFPZqtIuDaoc9bc9hwbDUtXaeUMdrTIRnuzxgi+DFotYhT99
LXbTJjbecbs/9Wn+eT/6fBu16KTpdA6ZyPnOCemkWmyYTI9llCXwNf1lnZFLrHxJpBZ9fECd/7u6
ZbdkdoI4f0M7WnX/ySXNB1myc3Tw5zbNBOrmBf7QwzTFoL/cou/+R7k2ae4FB28g57TQpSYuntRE
vGUI6NxXr6Vy5gDhuSjvMXDS34PWAIgobkYrX4uRfeG7Jk+8gAPeHKpgjtyWWrXYWYgj9WjmN0K5
yxrGOTLwsWSQ+SpEZetJgunRJQUy8DU2lhGMV5zWX7rAoPrPcXSr1Qc6KPOXu5p0C/6eGA2vikqu
zluYWCNspB0daGAKRtdrGtjCgisa1En1vYy3dNch5gUPQfxUky7dMMc0k17Btl6p5xnprxdqARH0
SbNSF5ks7Ve9O/NTt77tPJIaJKVPBsAp6WicXrY+y7f92qNOiVUb2o2Ff5zcWKu5YHmGk3PqMwtF
FxkWPN59/AVI6/Xj1La6oM0ln/0pQkBm3Ram7fpX8l094QqotCRQyATON459RMV68WCgV9h0Byuf
9vsb+36Cwj30ehYFpCot650sPslLA7Ey/6dG2E/AkooLUeZFLXsT30e7R9D0WSx6Rm2vrF6M8k43
8r/VALA8hNKi784EZ2Ja94yo2KJ0hMHbY8SGfEKr1q2l6c+V+2qlDkf+wLJd2hHroiUOz4UDxhfw
LbX8HzO7OuXPWB88VvEXQUneOMH+upLQD+qa3MVKX3ANe6S51Q/w/ULqHCH3GUQtsN/PVJ4JIvIP
aVhxLrc5I4SOujRaM9K38D6E0ichV38ILdFr0LBaAvMmmAf0UBDFRvEefSvDqwDuwNRbn9DSW1in
Lv94ZnBfEQ5wQIbn7p7PN8jkuC/ShPngFk/k8jcRN+vdDsgb16bnikvx4IsM8gq72+ZUcujU773n
DB+47LArSImB/BNKwx+rDKoxRHLAdRHoQ40K5mUPJXhfU7SumQPcYGkTRfrII94q+e3zFY2VicjC
9JZBJXyege1kCfAFrKo2ToyA75+8W2dn84FHJuFS10q/OJOa6Fn/AdVtI5lkm0EyPcLlz6+jqx+T
PoF2oGF4ekYtlktlBuKrPLzOGx9tYHZg+pY8s3yZq+kZarWttT+OC3pDRAhwss4AEz+thjqi2WLs
e+iR+54Q57EZBMWl2tw/mqrItEWY62MyriEeXXx3o/yBo/oFdnUePumw+K6ZL7j5VqN6s5yKH4h0
Mrl2c1NRivzacVEKDcg6FEV0y1JjG26AfCZxpkjy3HNiVXdowrVXbFUldlyVbZJ1DjBb8INhhy/y
rQI8TVyTrAW/IuiNMo/uE/1rwUllP7VIYi6HnlZkdXH8Vm1mIaQQi+pddFy0AHcWUWtX0cyr3T7D
564yTlkBFjAo++GYNUH0/N3QWoEYgzorWY/wS/ZsDhTVJXtzFqPXRbibRh8o5ssi6lLPzIxKQsOW
nFaLl/MCtq4tXhiPZre8x+2s83tsvK8A7Xb4d5YEm10rNvf1eU8nQkETFec6bFp6LDJcygyZt6Qu
iIC8Cb/s82xcdl1jEf2UqeazutcNtd5rz3gOl5Oistwi1KfxDl8OqX1XroOb8sRzjINUKN5BEALD
scYxecGwFkz/re0QFj6AooK3fc1uDO37+JnovsGkat47V9mNG/RIKkPmrtB/z8UC4EWTzKMSnPK0
fOJr33TTjSASRjcLZe6DEntHgQprDcFgaaInl44OWSsvdP48KMlF+H8Gl5cMFJsPfyiJbjAu7hxJ
I8z6uTNzamc/MJd7qaeF+p5+Xxx2KhItUxcFsoaKN3ZCr53Gr6hKlMT7JvOtFb0jlylnMeX17fia
AVeBz8iok+2gHRCM1Plfjv7RRMOQabP2ZMPcnJjfOGUgF/6Wwr3pA7l2wyEfplWwZe01QQY9iTog
bOOnXIGvdpXXb87gy0SZhQr7jLp6U+8L2gDQJxU8glGmhc76i9SHE/63Ga/z6wYf2IWatSthmy1p
sDgRgsv40xQS12jHYbU518PUw64OfbcChczAcE2ix2RkLIkt4NKVTjvdZ9aZj3BJDpb5bLJFnb5M
0XxzHxeY2CN1jLdhXDm9JUst3DLV49ZjwRaCASM+Nqz7Y5alMVd24F8epIUmsQiLpSFGVgQaBwYN
PU9BYkX23TWWF9hNdk/wEqeytku6loLNi4UHcCsEdUtYnJafGUDtTKr9skpzu+646BCVQFTPWy55
028Y4Ixn9kV7ucOpl4p4g/pYUz5P1xBePGehFTkzvyLcOSOfUXpiuah2U66C19pHUB5HiRfHBr/H
bgJ95lbigY7A6i5RWO6nSw0Cb38F8CG5KFl+vOZYAqVhXAtpdfxxoVaO8aPltyltGIcAud/yl2Vt
nIvCRVjCVhk+nQtIz3gOwdo5NCMfBu+jfVoGYIQUK9YbgBNN9hFEVurYCCKoQaxcTda/72zVcX7q
fbcEtpeup1LiNA6nTVujvtDqOmMYinDOmzZjAIun7ZniMPrlRvE5TiO1z51wEKD6zTEodAAcIdYc
Fwf8OGQMO5lVUR58LHSynoq/krT9nNjB3OQys3hApUwCV4dRlQY2CX++5kXG+3mwqDi1t1nQfxJf
fnHH8NsdxN7+LcIfLWrpPvvqpF8UKgFCoP++EiRfzCjA3a9hK1Gf9IG3N/VZCvZeSYUwQnsyj8AI
4fOk5h9P4ZL8lZPBck3hT/X9hWXShNgGfQ10k3sIaP6qqlyOmq7gDxk3I62ewzNQVkd1lpssWEyc
hhbY3CFL99jXPya9FJCzGhe5lPS+EIWpjiP9kFdwStzxWG1MtK6wazdUnjQey1UbikaTatqYo1UF
6psJYRG1GWPsbDuyWAD1Kx/XsDs2ObEU9EO78QX1ZSbe2Caj7b5iVQIFio1dmAeHri1YRIboE3ji
0/5DjympCrb5uPwtLHzxNEziuTmfhU9HEhi9IOdIb+C0+z3+pNGMR8qRS0nwPjsUfeSJuj5owqro
X23LaiJRxfoDJxzivs1tJ1IP9leBq0t+4Ld6qyhmq7sWAYJHgvcaNhM8fJGQmnbLV28g1OhbVrWw
XorMmuSKYYhc+BWnGlnFgEnt4Pd8f77+uT7K4N0waqTZNNP3xzLaGMcRNF2NQeJLQXtzl8F9krTB
A0nT15SoDpBuEOplX+g7xHaB34ZqPxd6bQ+Q2jNMyZjySJ0UpL78no3lxu57ansS7Hp+KDLSAELs
RIUAVhv5UMzYnjPEpaowbFx7Zkc4GbiRvYMSZeUzv95PYIZ18qLysCDDwDp40pFelqbYrKjVgRc3
k2mi6HlEVnC0+7sJVRkWvHL+XZ6BF4wdJ6fIDdrC8j+8nh2/8uC5XmYQZf/Wor818vmAhXq1Trjz
gulekmlKNnzaib26YBUg5kZQir36+q7X0zwG8X2R/XulxckE9sa3IlHnlRtEtlnKBkKL08m7OTqf
SxuNl6HxrMegiUB6OJ26rMOvfSS1/GFrE6T77Z+j73PHC55MAoFnCPN98IsYumdCMDJO9PqfNRMp
X15f6FYO6Y8zE6pw4QtuE9W+muzKmL1K+fOwEmusfbFIpkuJ2c/0tl0H6OHShyjCHo+jvChfyNze
PVSj7QvqPb8cEtth1KSlaCJbljxXK+Dev75S9KqAnMZ3orsXGr+FxG9P7Y3xgO+qGfhdZdWWX/v5
1doGjlbu6uSEVjzpBn0JqiBULhjVYISUWnrz/AIUjb8ewUDqW74vRSjTlPqw0Q3lNPVK3h0E2Qp/
5qJ8b8OLMBndpydDQ8F6iA8F6ZG0Kvlh5XhUK/ZSH/FIW9acOoOXeNq3YG5VYy2G4sa6XHDNwr9+
vNAbqWOLUbyFqtNQIUgIvUyIfCIaW+Fgv+75GtJoFKKnm2CfXhgMji1O0NJXjBWPX0YsikVlGPn5
6dBJxCPTgGUEzfjd8W4/3bRX0i+sBnp4ObbO6hyghU2b/Kc6Impx+fY9udBwioSKTSHkWMRdFH/L
Bwe+4veJg+CN97o1iGVRbkKUzlM488Ry/CZJAILVh6hCmgEdqR9A6MPnQj5X3qaEZiAY7keTg4xB
gDgI0Ef9yvq4jZ4aiuU40HHeYQbGHg2uubK/zpQOaz5XYnB3bV9QesngL/ykyEEKphLNofyxgI/4
kxhUX7/tcQvij2E1lLQ6mElIW7f5DwQ0qim9QkB79xAEk7iMwDHW5O50gZg4KrdOFDYjV0TcGZ/W
k6mJ+SgCajw4RvuCS+RyRyu9Z6PVczwncVBX5hwtb+LK/bcTFabSv2hAFOqh6UnFv86/HGvSIBtC
TNmQ3uh2PSM5AuMBwxmMiKBJ6MBKypT1mdGcy9osBRzuQ6HecD3vEkusSaoQWW1FsyduzxwMEP0U
n8ZPCAHThojRX6bSIZc0tNbZdLGWMU/Q+dHKoa+E1610e4Iqcz7JMIbPc114joD56Xj//cfB33w4
WJjGyPdiOy0S/+P3IXNrxwQ8T79lVZO915z/M309oG8mTljVrkQmWlbj5dclJZPLUzWxBTt4F5YU
tqmgVgUatmenTF77THGUmFdZZPr7VvcMZNDu3UpTJ9YuCcJkdx0qyQLJ2zyGrPWbIY97+ag01/Hj
gCDTEIMcKmzo4SuwcoyZS/dNodoKPayJqff+20oZcE4d+7bp4eXV5cwZabmDf/sr/y4jg2ZzO9/m
rwGaEbL15H8fUDXoA0+B4lxKtpMFQztRUHLJ92KlYMqFW684qwwt5u2+QWZYEyOzbYnYJg4HGQMu
Du1Nhqlym3kW8Mp+Ah8J7eCcnGiEdB1alowhtEuH3UxuZ6qDpjpWMWsb6lt5PwYKAAQg9xPUT1rp
sKv1vCgfA0mCmzH3BQ11kwDUZAta1AZb8Swn9ngX/SJxc2nd28nOidX93mheuj/ewNA34LuZg7IA
U3iKD3deM05xjIHcCTRyhro76VDTZGDhRHSHUep4yStnthrrK0xWCSW3tk9cjcM7u94MNKz2V8a2
gjpS6pEOJ1n1WwPwOb/Cwx/63RaLPEgfztRXiJnHhrkxfTpLinzEfIRCf06EBNiARuUJUumbMlAy
Zw5X3s9bjtEIN14ybpvXIVrmA1cGsmiyWh79e4zWPm77XPK0rb4OqlLCoas1KvaLLnz1dKXt3MK8
IM6YYWyv54kguqiQVoJdHMEz9I845Lft8qKWc/OnpW3NlQ9nQooYIP25Emr5hZCkVuHr+JmVu/Nt
ILyq69mn54hXYIUJzi0JNeM+yxUfrRSXFOOcKm4AuhUr2ux3rbgwoUPk/M6t/Bz/J1z0u8YfvCcq
S9KMkN/hX8+gtXlWJ3Wbcj+EBMDALFuV4xB3e3K6yohep6o6/cYUkthA9LiBiCViWfra6q4tUgsp
YSijYGTIzXTJEnr/ivya/Ki8nNF0/9eMBJruJeUB0oU9Ug9eX8dmuIJNbkNFpIYIzZ8hf4JnYNzf
WUWji9kedtZsuh7KUP4AI7oQ0ws4XGNRZw04V/CAFM2NYRJjkcJOG9SSqKcpQ5paFWmnCkHW3B51
Sc/OGIZ/TjuKfD6Dfgh2VXxgZ3c7zs/Xp2kQoBQeGCoXS/j714q73O98huZoCWlfUJp5PI60UJcu
OtYyk27b2TroxuicruWBjrsPdZ5F6cDT+0sIlEO3eA6wkfS2jVwuhZqCNEHHd0KO8vrSo+2jmQ+z
A7mGtnMfgKgElFSkSybBx/fck3wY+9jdzkYeYxSyQAJJ68cl+CKUGx81xFULTbemIj6vQ4je7KdP
Wn0OtVABwgBGuFJhVsjiNQo7N6N/HcD5f4YM2r2V29oaKGzBLKIv/vQ9MG5l/vE3OYKfXqM1UJUX
aqUyqUoOX4zG43i+yu4UF+JI+dcJj+juRVBhxunkZ/5GIwZDwljrPsP43dt77ht7ibHlkAM0qTlE
cd7pW94bYjmnJ/TBVu9/nI404b6X5aScDLvyuVuphSEsIPsoYIAlFTuAs7R5YkqvHL6ktzf7FG84
9GP8gVfvvgdwwRtBAjb5Mv/xokAErq8qBKlflTE/L/MhMlGKGKVYKiHpy9kbgbZzoj985DRLTdvq
bPC1t3bZ21v++K8w6eoFLOUctogGW+q7U8q5iY9ljfwJ2apvcKAgR2F78r6i/WuK6b8UadqRvuOh
ZNYwduafloXL6Xr0qH2pe7cau0+GMF/Bo/W5+E6L+JgqbEX64csbSUQCovdo/JXrWseGL5IpnHQu
YXq44PGR7csIcKhBthNaCfIn2ETaxlXb2MiwYxBudWRJzOBpf+Uobo6bdaWw36ETZfBIlpiViU5c
tupZa+4ZmCoRuCFUfYT93FxUEOlHusR9lC35UyUpEPSScwrICALE0L0bOh4Vjsq7d1CwL9FI4UHI
lSPU5Ut+TyrnKPQ5RELLwc3TfIF57NC8TkbusHBw+adpeSXV6wid63LRPFnfvFeH8TraYc7BAFCW
AfCtqEhQvfqZ8qupW9ps8+qGvB2LDUizMUwZAK+pDkkl1OqTaCQmE6hq2B7bNMEGCjYr4LcacCHN
9zRDt/Y8GqoVkxLmOdDGLtpjGqNWT6N1Nqbh3/qigLoaL1qYOmvOo6c2jajjR8HRqllQwA3FaSO6
eDpse1mJvrIDoRK6R7x8+yFKnFx8/gJD/2f0627BUyFu7G4PtiHv+rrkApB+PzVulhEAdTf1Ke5w
6Ts7UZE2+hlGUX5axeQwWdnZKCY4UBK/R3Hj3k9bevN3sE0EXgbVmkpPyyDLCs3ORJIRRgpb/zil
1Le9CLMQCrSWYHwZTM8sDtHjYEUCS0GOZMtR4H3ArsogBxSQb3Cj6P5q5r5KmhdFXqg2mxJy2iJe
SIKeBBoBdmmDy6ELtsybavBsHszAP+Iud0ZNYWVedAlAWy940KyA3S2INLj+l7fjFXlpdehJZ3jO
aqUzmOmkUhdUIIDpJ3kRynUKhgu41LqXFTs4pPKijwO95fWtXnEBeBI5mx+/aZHPebYwvjUzWImR
MhC/e0e1iVdPZMP65YVHEkYICNP2RmLqlU5oyse7L9vy2Yv5vmX4nbV/pkYbXheoNBuzI9JSy8tl
8c9vz/yghSI4pxDUbEssw5BsrpLmUkhgsSmTCfo9VGlxJ/cGl5/HX7NT4Cxxbi7A/wq0zFPH2bK+
qGZ+LP8o8li1JpXJlYIHaY2VlPde4wujYfHuVTJmzgEpONjSlXI7oplgtZ1BVvTnHgmLlwCNdR/3
kqwv2wwBbbnzokjHk4qE13MqgR2B8bIuervgOY3UDnQeiX7it1ipv5m//318IKaiso/Pa55odGp8
Y7WNKj17/bcZYvxIT7cNI0m/QGIAFvwKJvRKTYnr2vh79Yxpq0/xNNVDpn2J/oFhNq9DTbiDalgW
+w9asxUNxGaTo8XSjSAJfEOzXe5iYMdYz/7OA1aAMK//2qXfwa9qh8AONT6Mn0ldMPV/evpCS30x
1C4AcXuw32nGnHcPcnPEExM3RpkDspKjPt8lZGSv3ZSQHfml+sGKSZ2aheUxWoNBQuNFcC1KiDxN
fzgvmtxnZhZT0Dup/jH38Q5VjbU/+cQJqcZL0J+kIaB2pK7PsotU2hCPcyQt4hfCyroVaPlRowPJ
ybwLBC412kvwtyCZQOkPM5hriUkjmxlBvOf+4IP0vSglJhU5+1q2v6p6bC1xg1bPTNnovt43WEpW
KZjY57V9qgnMWy1INgymasS5IKUBbsm7BuNBwQH0qwd7wqBjRcO5XB76abCbGXK1AkpISlkClT6D
ic+1e1ZjWcjWaKA9WvCuwWCopsNZ/C4I882sWWeNyxlQ6Thv4AqtuLEkSCdh2TWOyuhZ1WOFZ/3w
3hHkYcuVXlEAy0yaLvSa43tBoL48Enjpqr7OJwlvM41otp2jR/C5JPfaoswCz/GYpf1l7d+4xjKg
h2xk8Kt4j29zyJfJKSHhqbZ959wcWJq/M7Pb/pZZhKcF/gtTXCWxpQouErnleDDcdaRxmwPKalgB
FFx6y0O4kDrdRhrb5z5TcAylYSXk5eveQTwN9QiAkabafHacEAdw0UbTDEYA6s49aNo5KcbRRfUN
xe5in5BDqaOkQfOEAaLCmcjj+oCibDcU8ldR8IW8QYyrLZNVB850n/OjPd74VIGhECfGNDzigdtB
6+iIO6zw+qefPLLtnX7V5kt1DMIC13h5CYx6n9GrTV/aWUOSoVQvHZysFIG7aqAHXP/eirbDFn8y
s/F42SbGaoAVwBr2w5mnpVGD3kKAXDn5kCFvfIrtdsyZDozmpty2TnlE3MwC3PC8/+rrH5d9y/lw
M2WOQQJ9KAd5RdblFD1yAM3ej9+3HGp+EWzUF5qpR6elPZiHMh6DZTjyP9U742G/l4qAndDMFMQP
cSn0KzEL0onkjyjokCOKLglU5o5VJ/rJfLjHuf4TfXu2FykV1Ehn7F+miTtB4rNhR3sXGFbylG5/
hwFu43yvbiI/56vigyEPxWYMR4M8N6KXh4PmEv4J4d17dBFOGf7YhN1Yc3zTPaoWJIRd5rxjkBwM
P9G2gXmm1dxZxscgDGFZzZn+hHqiRMEai6ntqeoaW8wwKm1Z58O2ZmzNvTeZn2CYsjveRP5TWHVP
8R+VcPyDl//rQpVtO2pBhxEkOQhzdXDpsF9YJAa88zHVYc4w6I66Pluod//pfNouyLyjHtbL9fWE
+mj7Ffp9STu3cvfAh880jpiYWLdUwE6X2l5UGgJXhDONi1k2htjqwk4HDysQqaQiFiN4z9SF2bxN
L4Y02N9YDFY7I21o7SOl16H5U00L5U8N13KVGMdAg1siHuggo463sHhXF8bCvw7/Nma+hVedXcz5
b6543X9b10MjqZEGi2XEF1+GKr2nKGEynJlB1Nixv60vPJe1wNhs6e1RwGpkgC+NsjpozJy07NvG
EXo9ByPLI8i7x4/T+EoCneh1Lny4QCEX3jOhvv4JdNI+ONVE3CyEJK4jbyeY38p59EuHBs/619Dz
CcwfRj3X6SnFVX/NxYzKiSbspertUR5Xs2AqT509c1GnHbw6tzUUHDKfTpl6nmEak3Bd3LJPXtwp
Zk2gxZPXw5GPrY9z0MPS0y+Ojx3cCbFEUFLJ+44uRHCtsMJNDHsOyR43S6DWm73SCl/oRdQHb19P
Mnzipk0pPkGBa+c27f/VXcXRA09UUu0XtBGcX8I5ae+uTxsmc3DLz9XdCfK8OdY4S3iKGczvuUBW
AYyeQKeifVxeI4Z1aFQ0S4lqA1mKo1nGK1+XNOK0DttKaMf5Ezj31RgjnGj2uLhaPWWSwvz/ar+j
GU3dL+eJP1CPHa5ppegCRmp+RcPbYj2T9CjDTUy/6XUdvWFySeSmB368lPDizwXXDqAI1baP3mKV
zDEkY/WZqNUbhirDp4M6ueKkMxNzISMTg9txHH9qFB0o6nn7sjHAJMsnQKGMfClOfc2AiMJsgYmR
rUD9rAp1NnnPnAn+L6YuB+vEOzDht9GuuUC6tMQvahHJunbWAfmOiuiUhajp2OZSCNO90v99Tw+R
tUHydlE+kC6xyrHhVmBvotRgMMLdOwtvi9YbS7pGpabZmBTDC4hLqxq16MC1JCgMMWO2hLBiuy1p
EdB0Zn1b/3yxyj3JiCHuGlS/kUK8Ec5F8JcvKsOU8N6jAgjZK8aIorvYTnce4tPRaGy9+nE48HJa
bBnZ+UU5/JlnAciHmGDPN0jSVq+FAAoDv7RCQJ7KajglgoEgEoEO028aHpFa/eUvNGdw7s6SYDyg
1kT93uQ/5UycRa9Up/k0SsWiY81L0bRQ6buLnTvXf/y4VJfd2wnRNUHSO6vocanlrp3BAQ1YfV3G
HL5XHTrwlaTFI87Sp7++fFZVO1jWDuOfp15/9nOfgFGVJgOmouF455pIXmhQeMGnk/5ZgTeUDnR7
LM41rfoq4Mvuh2q3Qa3xkC5lQyaXuSUTfD9pti6bEUPmJWX+OUunRH3ptUnM4oweE3/peuFR/ylp
nSfBR+/+Pi5kGh8xt1ymtleuNWndW6po+MPuuoJfBDRAcMrvYdMFIW7v5J4E2oIj6knNo4j1elDI
bPOWQcnDX8aj1xicEIBeN2vN/fh4PF7LgYfpLOdjRMWjwQuoZELAY1ApU4gNl+3I6xrYII5JyEDi
hhRspHpRz2dktshWc2iDadGgt0PG0PQba4KTEOzM7r3Gs4dUxRPIhg56bg58XVTrFCleyRqcrEQN
Q3eiJdD4Ws2OnNk/FmHv7N4AhBy4i0DEhpyuuf5vbofevGGRcL8O2/9w2y+6TUIX2i27b0bwM48Z
sGDSO2m19eP7BVm6DLfNDOiF/NNd0rVxGq/jv7Io5OEVvcvSUfriZQZ5+8hBfOXIFGDxarK/l3CV
poxeM+KK/u3ltHpIRpVU4KfbMxSBtV7Nzn7cAIOedVLTdWbhLmLKmhTrEklR6WnkI+gs31KU+29C
xexSu6uhHitz2xbZ+cTqFtvD7SRzAng3dYv11RDkvBlHrHzc+e87RmpM4ghGtpQfqLVIjeXeJSrh
wbeyZzfjvsp2hTyzIOJgF6UF5PbAtMp0b3ilrgBeYyxQlX6gxThz6DrIu3v5xPGpevetonJBNpfN
xASuccyBTZ8hbYpO17j3giE5ebbN/xwZHHekLyk+8XtpH/uOpR4e3oDt2kJkOFJVnvc1eqzc4fwB
0lkDD4pdYKmEIPJSpRGLZABrJdisyEoA9mK1ji8q8ays0FxCuzZB6ShcqDKCtZFqN58RJmhMpbqW
3SWBmRrgqxPrIyID5KjmjbTNj/8HknongXzlFjKnO4ozKjULQakBUBGeCJ3HXEX1UCXiUDY3SQVW
Ua3BGa4V7gILVFH0DlF1pFGUuj4yXETICyDGI87bLo+edD4bc+EvC35I8rI3n9nxyC4q+FQ+8zd1
DjGw/K3RRrggus0rYSVI9feKVDb3cxKLD/FYsqZf00xQGOQSuK49bURdpZQ+Aqa+w72Uzc4HfOzZ
Gt6ekOVmeUmD6bFw369xHNquumpFhhSe4SSc90XgdV4HOId6+OhBFYtG4yFBFjZwUtbBT79I6TpR
g+hqYsdJM+acvPfMzeRJyo7bZeqA3c25r2TfKs5+DdMOo9oB6wXHmQV3z8gqA1KWquMZkcyXnuoW
rysTIGX1xXmGmkdffO0kI9ZMGfTU4QlZeEMWpIx6Smcn/mzl1JKQD1IgP7kQoS6JfH3NSOsuz5QS
rsfZx/VYGlrXxOf7K2NsiVPUUmdthkYK08y3IF1j8kMxtCh5LQi/kF5UTRPIQBkQJnFbO2UFrrFr
ri8allbd5L36SlCGqzWGyFpmHKRqbRzLyMymyOVs+LcFCtEnOvg7H4kuiofoQsVupnRQEPcc5D/4
9MQmuX4pMjxoJJ2xOyKameq2T3xK8eVo0nUS2TXzKDRkR0Bvk7b6GI6V8Wvru2Ld4FtrW6UxFmNE
BaeYfU3xkM+g8KG1iepp6266flRHy792XlvSyLvZMHX4hOQ4HrAY421q9fAXZ2MZ4IbA15pgZiZk
JKmWgr/d/DuPss5tTznTHr8gK6pOJc9psJ/+sgFavyXFZQlPCfWzdtfG/gLJTyt+VT3J0BePtD9L
yGNDTvPqnRBABnM2Vyf8Dit7q9G/ngmcpVKjHtnAmdNE8rwxhdfluU9PQtkNByP20hA7HjajY/I5
Z8DZxhI4mUp4NaLk0Utf94DCCRIaN5QgO3pQH9gRQlOsc6VS6MnBLRXFn0Lg7Kz/bfs1tXLZXDr9
wAaQqi19GQ+SJ618UuLWNYqvYaKq1OSHRvJuD8t6O4lVS/O51nx3WsLUfhSXb8R9mvg8FaF2h2RW
SL5EJPV97ntEvjmXVHyXscIHxGytLhVpE7duMEC2moxKBS6GVUZgCnEMK2V+ORyCSlu1rHTPb5jF
eaJbPVvOavj7H9xVc4bO0CoiIa2IIQnOnyz3e5n//AzHt+4iLyGypmYLk1JOc4/07Za9l7tYc9Hv
Kx/iAFxH3sRsLsd12Np7H28QS7de9ofUtz4OUuy8+FilzJRVJ56l/9mZeg+hPCCpRGjhw2/cUP5R
yaey7m9TFr5jVygv+7GXw/BXfQC5oC1OYUJdy24N++4cuUXHDRc3zwDJJ/KOQyhajOZBEi90futk
+0seo86XetOo43aRYAZAjaRV6wGo73frO3QKXCcPGdTFsUATm+9Agyj7O69LeZd6T/yZyF1zozgt
LnmgQlhRiUtgbuMsG3LiLndhIBdvySK7GkNkQ8WidhmW6lbt1bTj/Di/5tvnstdF2x4BTxlSvUOP
GASRZ9ErfhD+NuUBxqUVE/4lEmdBedNHvkDWW6j4wPUDU1y0zyny4F2OVGbjfr8Cl7LkgeXZD8gU
V2n7cE+Inq9/bzTVuxA45oWzi9Q92StY4lg8VoC32oKlAKd3DYNfv5OKfDPRqXlT37sdV18+j8YK
oUCLg6O8C2Spy5qvDdJIKUS29tAcI6NvbDJc62S6wSZNw3IIJZ4RV9jO1DwAi6XBm+N9+MVDjMip
mCdl79z5EoMRMwdcf+RVkzcxOMMMqjW1nUoA5m7i+31bVVfNP2JCVCi0idv2E89nJ7e3qcI1tydc
kFhi+U2ASSv0QQFaPLn5o/7X4MO4A9qBLoH7kLkJdS/UUDPWgMC95yTOcE/zStnz/82qATNrEcyH
yef0JO8RC0kTKH/f3d2392bQFmCjEoJvU2xZI4kMo+igCA1k3zhFmI6na5TpdSFpxbN5qLY/F2zc
q6+I843hfRfNRxmKdR8ieMI7pE8G9hys8Avst1kbxhw2fxVSJ83CZckc1D9ItRUkMmULgtNap8t0
WYyVKg/D78Q9nwiIPNVzql73N6mfHxw4wIBeSrR6wncrIil/T+u1Yv/oYhFMbEyrUdRQGaQGnkXc
I0YR8pKsZtpnzfRDTc6OxVDNhTeXlbm7HIUp73vkmfvkHYuT3rgnQ3CILQ63EVakwmjeQzXYU++h
sF0DNX2mTq6wcbJg43GJWDXb5xE8QIFzQk8IcPkd2kzluqZpNeB72fhfU9IPIl0NnLMN+woQk3qA
QEDgFa1irTmgHzTEzpo+O92y5YbXRxaboongfnIisB2K51HxEigu0yl4miWyy+LtbFU2QND2lwbf
rvzcWdowxHXeJO7Ctl3vBTUGQAgnqzqbMKkU7EVFMw4gSh3eZOhF3Of+lUIRbfwBthbVBhNmsT4a
klqrNBI6oqQUO14NICQy4ekeFLjKcRrVd7FV/Nsbku0sxfb5jLt+kQR/uA3eHkOAIr388LxJC+2m
8wxZ7SZvp2vNBq8CBq5/slOHE0Bgn+LyjRAyMfNiROiASexmKQ5VmY2nsqqEUzgnk8iDZHgJNhIB
vViWKGva3U2GuJ8vJqd0gHs5hCNdJI6fbhJG3lFmgoXKE5GqdxBRe+GUJ/F5+/m56ZpCbps3U84K
hKbx7IxTf+wye2GcsrPY8gL1ldPNcSVwgAtJDNLOymAU3RqfZauF9C36dz26DVphVR5Kx8vl8JxQ
8y0U37yH9QXgsOib1a5GrBvRNem2knY2gpZ8CPrO9z6HxlN/IrB9RBodNnQA1XTwE5LOA0JiY9lr
Q9XKNS0yAvwPlWhfJxo08OkTfKnZbUBjY1Jwwchv8HD8pMyfR0T7BoI/mHSGGcNG2lnIKjmKdfTW
xu07FX6RSeBeOgkSpprX97E3LYMvMtu93V0ikWw0pLn0mlzcYWdlKi6Ao65PHwYAVe8//SQOyB7p
tygVu3fMlL+n564xdznZ0B3H2pHO86j0w59VMbjJhy6DFBtfZsleou5gBRimsSOFC+/QVrVP3Ckm
sc8Zt91vHaSaE5xCIINyiymNxP21Zzvu++dbfVkQzCGZG7ZniNn5WxYvx1+7bFhCjHrYGx3FLjyT
Wq9lcpV6Zsq60eDfDvyq9RI3ckj7ay1T1kCcZLU79U/c/Q4i6v96XXqskMxzS2XatF1apIMKdd/t
ucwG4+I5HrDlKtRSXOfkX9wj5bh3wjJ7LG8Rs/AwzEZ6/T56E1WNfnu9osjdk3yNxxJU4RAEU6DG
Fcd3wOVM/nHIzlr7T6qbiO7DUBGAdl1SEPDj/DgvLwFmSldpYzuecFlr5nrLyBLbsMDiuk1C/M2+
8qorxrQBHkvqggs/jLf3GzRgv49ZTqzprhuZEyfUqA12oQBeeCLYHDke1ubDTzrPAKhlZFw1QK9V
O7IUtTTvoq0Tnbx9AEeeGHaG0N8P+h8VKRjXrKp2rJTB70PDdW40c4z/nNop15lnp/ElkG47dLoC
xDp5OtlVArbGZn8aIVvbtiFHGXFBGGg81IHL4ONKSriz0bS7khwLohaQwhZ3PUYPPzjukggx1wfr
5vGE4xDFJ0+DM+Ah7OH5a5iNHXeKIm1hUW/yuB3yHtx7ml73ZmRftSRUNwwJ8sd0cbzsRI76S1xe
qrMH3TkZO8FZkDadQD6Ny6ENilsOaptQD5sVnDTaxrRdEn3eYvUBbC3kfMMY6s3JyCYZBeqDPinh
TFNmWT6eRXiMvneZG/MY6LdwIlzk4Ea4ILMNqqGF43Ygp0AViffFe7yvH+Wu+XiNFVobe0wnIWLf
t6DQ0VXvcwXJxmm3OIESIdCvRKXZf+TAKbcWA8Ucdn2Vu5EVMMym9626VN0GA4IXfkBGa/Zn2XFY
Y9pPfUZW0PK7aMj3MgdHvtxoJ0ImQYZh4ozOfXxVILxy4Y6J9EMZDF1qaoevQkMXQw+LIsyE179Q
+3Tl5zwZZ0ijZmP/OVJNPM7nGsQJqwujfvRPC568iwtYhePrJ2uOaiELPJdLMzhNilbg8Sbn18gJ
G8359Db9MEXbRQxoZsHLy439YXXIAORzZRaPzA5LF+puJi/D55XISRn5UoxNY+cZLkI7jePWsedH
oM8wWYD172riGpDoaM7HgomP7OuiZjX5Q3sqzBKJ4MuXY3BNhs6L8dlq/siLPm7nTWu9roWSTiEY
pK0VLrzI+wWST+ZuJVVibg+SZFrpPS3RHDvLjp4h7waRGTxaG0sSkYPSbAG15v5u+V+E9u8mwLhh
hpON14UmhyjFnmg9gWt+1iqlLPKmWPPuDVX1FAjeQXPq3ZSG4sxLvM+oZhxcI9eC+nfx6EgcBTBw
tRTxtmAFXfMRW/w30M2tjw6PN1fz2HzG7Ucx72JwWpzlGptbBCi9ApMUfsGJVa5vn1k6ulaRCAX3
ANH/4Dn5bKitYgV9Z4DheBo/SUfYfEEitLDHs/7XAlui2MlNAb2veWcYs5q9fZTRnYqUxISD6nG6
gJQSnQchIx6aqNiJOR1kYDUMByFM1d8bFCkJrG64oWbTvzbrxGsvI7ATUB6+Yh6GSrI48437gyDv
oxvgaRUHYmdw1biq8VHxU6q00yB8lmgOOE6G1rXmcGtJdVdq4uLKHlqkjnwPSUm9zqrNXxYZhZGb
BM/xZl8L8QST3bmh+V0Fu3TucwOXxhlXnYUSvet67S4CuIJlr0n97eP4hODz3Q4dpz/V9LOuWWLd
+Tbxopra77TLBIIP6Ib7jqhA3yly/RVVSnhZIzSx3P6nT5Km+Ju+qNz3zUsowuKItKasuVaNGsTT
zNKOUPDA8d+z3QnIqoKGKivvfs0kWOgiyTcexZGF8kJovIP0XwdBSB12VoFcBCQIeWKuPEQ68gNV
bd4LitiHkdDcByZro+FPyMvYr5FX364CFKsM+Art9nsBCX1UPeAhVr2Qx4AbgEbGuo00XI7NIUo7
H88v5oNodqKRIFNsMjBdyEZSokbj4rYjvmweNlgkvI7P6b8dCLsSHqfBIQhKLdQ5QFf1VRVsxikd
oVTSjh0OlMNuvFDiA0xroe3JJiF7miMsfyBciexJTqDX17o5jibYbtwr2gGDtVOduO1/czE/x+Zx
2JZCLAiAzmUwSAr/QPcfJ90WgeIuNpShwI98paT7skcBIUeLkgXgROcW2yqnL1axWjbbobnv6cjC
PWEtH0D4uJPX+buSDcaooInJPzMfiSahv7syddizJsrGSiqCZcfTPve068uLULSPwWK+GWyhXpOB
m+tlufBpxcKrcCpBPiov5d0LXE/vtnTNF+womlzlKadbDJN/r7s75y6bu19tVs9C9wl/zDd9qlH+
FKhRSqArq+ISXUWdoO1V9B8Z7p4ELAehWhb7HyZBHtgRujV8Uq2b8p46CdacZqpVrJVIBfNicU8s
ZRHBRRNVWsK6/mr9H79bu+Ffbph0vHQ7TnXf02rUAw6mk/vB6+SrlYfqFrqLHuBg//VYQcq5TSuU
jFGbBBndi/5hsONg5XtzBycIZhOm6C0A9tHVrwmeGG6rbIRUZSGo1eFoo01IgcdUAPmsPEuJszhU
iTo6JcyBewu2uNEph/Q1R5mWD49nCoULUGEP15vZKfihjEykk8QcQbRkh4xkb6gfL2EP3OpPfICJ
u4uyExnsxahd+8cx5ZW212fdYGkX5DkklOOG2PCfQh86Hr6GzCwzEQYrl1MmDp2DN2V7A5ub3VJx
LENVoF2EIy/tu1BWBJzWQrvtGV/es+WRpNNKi670gfvVggv4wdhz4zRb4+yevEUiL3eXxcyd6EKG
cStd4yY8t4vauOdadUOvbgf4KupNctzpoyCjeJj2I4odHW4KUGzo5j7MIkgkJhLmdFDbzD180I8Z
op309udO/iXWyCtGZ4zqznNRW9uH9M5aK8JbMHV1tUyQDpEwc7KlZAiMBSLiJjkfF3CJjir1sJNZ
WlwZbAApcqPTTDoUOx3RzOCz0lVkEipru361DsCvMP0C/UB7t3OWF4KuiOqueGmoxGDEw0Y9yIeu
jAWTFQnNkT8zuc8POFLcQVFmXkHKyTPY05Sz4W70MtSSyEIpXaas6kc3UFMLnPpXEpWQl26TcntY
VukwM9HEw4R9CRdnvaHlHOtHdKXmQJyVygvaBmuj+URpHrWnlFrt94o9spKQMSt8THLttiwJB/M3
h7XgrDWEmccSrk9jCIBNI+8JK8Dvlj8PbJVlRGT8nxQurptEssIl6J3c8z5h6aDp9YFwQdVl+Ha4
D1IPx+PTXG+WXseVFiSm3LQXV1ppNrFRk2L5eDrf3xx1APP42+XGMvE6ifAnFzSQgNSDBhI7WBRJ
cnJjRUD8cISMw2o58ChF9mVPfS44l9tfDzEfk3R+dtFvCd1Yzzd8wIcUhJpi95m1jGECbEgdsCbo
YgP7P6inXXXYRJDb/aCX1hyxGNqGX2zjxznrCpiM3bUsAtZ5mBrOggCpiKb+KwOZrYC8LIFyhTwP
9GhS1eQ99X/ZtyWkNr1tetx64b7ef4+Mn8mpiILMYF32t1KLNtRJfHnm/9Uf+cyDcXYvZ+oaRZhW
BAXJBzIe8pYIxxqXVR+9ZPJAXKoQZiHJY7R3LIpuwAdqLut9kQbHzAWe8zaUqBKD1ViN8ymr5OdR
EUABGQjo7QSfcfn+U0v768a7yh+TboGJlCLFAEWsT7+VOxPBiu+OZOawPJLkk5PCJR1KQT4NQIpZ
fRqMYbl1+wP/kdFTEZTJ9qFtV1Bn9rEEzDQWwSmBbhSd1IAjQf/hILbAeV7rHf6IW5gyehYmwRUf
HMwQj1VR1nlIroDPcsKbHdNvRlurHovN8mGibEKgJPWThksOaKZ2284iWWiwWbFOGoLMDo9nTITb
LsjNsldeX2iA+6HVfvSJd+BmyMSLPocy7AobOura4OSruvTpQpxAh/b9sBrBqYJTfg7VPFPkT+1G
BsiPC/9OB66bjssmpeOtSmcjr+xixSFiPNJO+1MGx1CNDfF7KC+jbM7gF+QV/LwI7cxzrzH/+8Xm
OcLMK5c/45g6wQcHXNtXKp2f6A7gqoh9i4S1OPYBEvnRNvGzuxSmK3dqQMW2myemwDiQ4SyF+IhF
6jhTFVxP9B/jn6k7AxHe7/Jd++kuI49HMa1OdkN4BWWbzqMs8K1f8thJtbijTRsfGe2V/YIAOd4I
Sy9xtdqHVySHrtnVfFQ+jmp1xmcvO2Ujn+zWmU8iUwodCLIEZen9xwb41BrFt2dZF2A/iIQV3hUj
e2SGb8nGCcDhfhe9r79FimkHgd6WqxartKn0G9m0zD6bW/RtbA1fQxHYpHEoyDhYxSDNY/n1FvrU
dxrtRZU4xYKuHBptMsEwA2MZppnkEiMDQgeZdKDXvluwiLD1qFXG2Ghat7SFQ2ME2ifuO/u24VTD
uH/Ei203ncSfCW083gzWbBmQ/4dmgK+W/rE3gyvgPU1Lebc4RL6IfG2Ulu/2QwARD3K0xPC30fvB
5JvwmQaxE38LHhzZYFDl1gvZbZiyD/HIlCumnX4GyjATI9JAmc6sKkZvBtGWpOmbmZeEQFUpDpaQ
88NuMBzAdfIz22yFa14iJOmerRRoMXN5hW2QRJFgSD+0ZyNHayx7wNG2/yOe3GMO3nwi8uXRzJav
NAJmy3KDy/VANcvmORJCH9q7wkaEn6uWhKKQ8aI6GYTcl+XI6RfnMp2C4zXaUdJ3LcaxM1pula+x
po0JNfGTN+wh3hlDg/bdVsYcEowGEZ1ao73nQvIF1pCmn2ily5I+T38XZ6e35hysRdZosfxLobUP
0B9obDLqMoLVl8Fnw3W1L5DWJdWPOIwpAmSnp2jSHMs193SZUKTx1fMS0Vr2+m89WJdInvFpD4w8
bx2K9XH/07Pqx500aGh8C9IrdIwvjHo8FEJ5U7aQVYB+KianpaTB+Kd8adBTKtPjQoZ6TijK5u5y
qu41kkm+xMr+CtzmnLY8nDq8/KDQIt8A2fpy1VOrvaHfi3QDAgmcdK2lJ2K5dhmzxoh9yyMtZ14h
wYzlFYCgq/oHsv7pryrYZcLOlkP8pxBMjOizkNivWZr+PmyqlHEbajUP8PilLSOJ9ql/fegVWhR7
0EXl9S4x8cRWSYXSm+7D6Mm05AXmmPTaxHPZLHlFxhSj+r4FXCjY3D1szetZJJZIu0JBPRTrXl7I
hlRCAjUp+j8PIBLG8jqH5kZJXGZRupb9UE8grlIh2HE2VSSLmVaDDcFpEYDZUs2Ckzxk0q2Ui5IL
bXC2Fx3spTIULc6wKgmbT+haHp+cjBkhzILN0Y1Gh59VwPj76Wg5/EdX/tp2e17r/ovvOrr95aqD
YV8W+KYEZzMBx0O01MyblXiiZ9qpEbytUPeDlrGQM88Ro/mwmo8sEs4vdzJngnmkOSEV/GEnnOEI
Of4Wwqjc52jICkKnlnNuVi9J+nYW+VlqzaGHSZPhGb9ASiml77okYxEMQdRQXBO2ztqyX3jUF3VO
POGFfFjnm/2E4YTxmabyrMuzMO8O7W46pscED7kuiChrRdVCzpPLiF28XnRsuzzcowjkSeXBT/BV
HXgNBfmhDHFt+VSS2YZQInYYQPvSbeZBmNidzep2/mC79Rau3vjKq82wZkH9ietxzgSGCUt9eBJ2
wA/lfUh0ZyTpCMLs5O3qJ63Oq62O3JSzcNuW7LE19L02z1M5SbwsLRg3U1zgGPWpDUKd+IvzdZPd
1bSzSReAI7x9iZLT8eLZ1xj6r34t6CPFGQGQcGXY0ttRekgn/b8086fVYg6l4GKIP0T2UyeuqRGb
Is/JDUcaMzNehmts8Nw4HadIhw7hygBXgHWXvDwqgb3YXCMc1/NtevYNN2bRhuj2EI4oUCqq9kc5
voSmO9EgWSAHrwSqDhC3EbynNT/YIzAd5mVGRRi6Vf1M926RD5KE5k+JhGz3cYNkfT2HgBENvXnh
3VwMToC5kPmes7z7UFf7tMhUzSoMcnPJzjzeAn/i44QhOHu0cYbdDAEB9qdmzkzeK8P/698/Mgo5
+G90bCMwXStO6CUtNlsBZkwJd7XQiIubjEG9asxiadkoyerWBsfa2YL7Yed1IT6I0xfPKY0zuqJK
a+LFHeexyTRBxld8eShYtjY7ezA730zFWQvo3KAZOHx7jtvS3xVvBZmjflV+CxrXjIvzskU/9BQn
a/agjUda2npRo5uH1EpVPfAvq3bs00phL5asdgE9Y4eOzcM2/0u0xfr5gL17cSCOPazJyBjqVMgp
usBDeeE4O7THIsdtWQCfLcjyfFjJcb2Zj7AnfbCgP7FtS1PG036HwDTloy53r3pt5+0N7eYTT6yd
1L9ZU4gca/3+jXo0+3v0+Qxp+ekXo+GMguEBCiSmsn7JIbmr9Ndt21ggCwDaW60Xtzj/+bRA4Xhv
UAJIQ+y28UkWKMF+HIkfqnJxQLRdJtq4bSlHVKaoPTRvamCgg7Z6A7PDsO3L3cMEMumGr4nwUaTi
8CgxXjTC34IPFqcGUAiJLMyJ1z8FNsKUWYUFaieLkqapY9QUL7zTECALoJK9EgKTScs1zouevNzE
mF5PQgSSLK4GUhxtxNA2KCpVX5gt1+Y4AQe02f4aiNC+v4JHo2/LGWD/X6nK7S2WmUAEGK9XHjtY
AUVjDXA3nM784ra3fGZHgNMVrpTHZhbvCxdzA+zVoUX4Bu46j2UqM3YiRY9vmx2nea0rubdyuf/J
D6YecbCfWg9C3sRwrCaXLjLxHEl+npAysSrdy/FrD58nSTQpfuosKPJag3XI4PwSQXcdzDgl3AeI
eBk+VxOP0h1Ro5ZkddF+A7Gvn0eXBFLTv42xxpbbtgb6lmKwmRuKrIm5YZ2bJ1EdMqX4rF7qX9WV
kcbXianPe6/wCR5frzAxZU5KHp7D2sf3oCYBeaBFBIMxBkrQ4rHFIiCaKDllZnFYhbqnVDbY8xoo
cp37Gh1qs9AFjvzuzZ0MIJfbEPeh0DLI0P3reQIjIBcgaC9MAlPt9z1uD9MxBI7deOtOJanGHbOE
vgwjsRApQiqyXZMSz60cEVlFt0Kzia7MvjpBOcV5pRR9FGd05/zUqS23UY4zktp1izNCgPdF5sZe
gRIHhCdmP0JOJSPNIHJ4FKCxO99NgKfJeLgUaXPjIWmsAKMjHa7VQ6WQunyQYWkY2f61HSkSNVBy
GCjfym+Vez1StmspR73zvwX0E8S+POxB9G1ocb71T0JxoZy9gw5b8d4Ndd47Dl4+XXrejlEkUTVN
AyExIEL67vEDUiQYkTJTnSVmSHY0YRw2/6LO1SAEe/e+I0R41zL8uJJc90thC9mdIpZDB3onloZ2
WDDJbQCNHGFEETyGf8ifZoIFo01TF0YJdaVHQjHlrQ2hPDHoKFPjwZobumLUf6+nKb6A6HEzoRoq
t8it3IVZFChrHquo580zvmWjueQrztNvXDU0ZLezMj4c0lfDjfEp0GwuyHOLnAKo9f4KYJiKRD9v
zBJVSzejid5Woo0lkoXwAEnazsz77LXQ1OLzOkx/ErfuPnpHCPLz385NY8iL+cuG/f4oshnoW4O6
EaTOtxv2aznGcm0jiYWf9ETnQNQzcEEKSRYIIF4I7qY8KCiw0f/Z+AGm/Nmxg6v17jTdfIvTJdQ6
lH7vUcx8LrhhkOXf6PKC06MkXPk1RmuzZf1kSr6Ui6yL9OwK9Yz/VTFreHvxPeuARWkPEky33xw9
hEzCWOU78u6GW0sdD492Jcgk4Z29SaP8l441/VL4l4G/jGL5VoqaplS13RB8T726IqYAToPv49g/
iAKvzPqjYYCBiycWnI62BE2me4Tbsg9QbzXHqOIguRDe9KyUB2Q2sASJemwbCcW1e3upY7mP7zaL
HzNB+Rf3yG88VDPykASkVAt5ONBP7VQBEzflloqAf9hPbUDdffNzaz4jCJBrgcYaArw5OJl0XCSb
Fn0VhW/FIyMNQPcqWjegMDt1mcGdiSP70kArEPly47IOojmZb0FkuKo8hAgDbLTAZ5bKs3rWAohM
X/NTI3AAa+SUGj/CS/3jFJXh2023Ke5oN+1XMj2spwcYUH4SpvxyCqV40LzB8OIgiuNHtYSdUrMm
zl9MPNNI6JDjYzDVF34eJdzHp3UQ3MqNayfv8G3fBIBEBMPg1RTaLbJN1G4oKNIdiU9ko/sfabII
I0/bVC788/+3V6DTx8xE/gV9qJ+1uDRhNUTSxhAqqVMoPoIkEyoglxLZ/umKIIRi845ZCNqjfoQ1
IrRpdutwuYeYdau2UM3bPj9BlGuRgA1BIANrzgzWeG0aSAWQG2eVjBpzjrUSQKOHqhAg8A1YygO1
nRUuMVQbK6USI4CgtRctoV74RhG4KZX3027cToLRfBWhLB55fySwQ10hRsXEvK2m/iJ1FdxzzbWb
7v+uRIbD/fkQd5hoGVjN9pSglpnFLELzz2s3t5mH5nb3p7nL91jFCJfVLEZlJLGn/P8Y+Xl1I4FP
nwyc4wdA0oaphA1JlHIY7Lyx6cNNpFz5ueJWGJ3I3Sv9+gUFZT2+RJdBVDISTjLfqwiZjC9PVj56
GswoQjpVpUD8xtt+73ntuWGsSbYn5/kxd3sO71GsBiJ8DRQArcMLbrY+j751qNNey0EeXVVjh4Np
jAaQtiDANjYnbWUbyuE5n6SBd+p9XqoFpp+M7KKaMJOlwTr2dNwp56DmkjMQCXzgaIW2SiWOgVfW
AJCgoupe9/JAANiLff5OzznQb8frtJKiMZT7dIfd6YWUREVjYA3cqPJZDWt3cnKGepUi2AWfLG2X
R+duqZ9Bz7hBlF0riDIl89ET6tPZmCzPnXr9ua0DOTpjBrYaXIZrE1z369LDJ03QmCrvf3JxOHzs
dqiN1F2KgWlzJ2q0UaVCiqUMrml8IMDQkDFw3ecVC/eVOx7vaI8EEXCr9opmBsHTcGJtqEgTAsgM
jgM0/iZrkmov/p7akyqdYIRZOT+uwcDoXHYD6Y8Pzqq5kPPrM6P3OkzBEO5h3xR06SP2f//vgJS4
90FssCC+4Cl5UyAbUVbhGxCK5LzEKULnO96hL1ZI8Gs7s0ZG1+f1TVvfuSNpslRb9R8yTkHxV9ZN
yPj2yADE8Vbzc0bqu6jeGTbZlpZ9G8rHOD3/StSCyvcrJD8qPujvkZXdaQ7jO9glLSGdAoDVBoz8
Tz38Hpc9PPHncCJ3FNcF/yJPtd3gWQYIuo2NGJSGr/OulnzmZVy+6r/olNkeiNNRxACQbYdRqbN7
Y1uNygxn6jsVdzUGkho7K++e2IxzjoYdyKhpjAYq/TJTbzGkNeX+fIq2ko81iU5UmRwhN5g8vN7u
0ktL4oie6JMIYJFdbI/FzRFTFA31q8WAXksjXWUteFaaTyJfhnCiMctF485n1TiwkLU4fiju+8hr
HfN4pTV+5NfUrQEfQGZOw89W3lpZ4PNU+8AW7DiaGknSCGaJEtxIpUerKVCImeqhRDGzIHwPd6lF
HHUN0rfGnCpE5EsxwI59krjrX0lXHxZ2tZG+omQzYTyx6NF3See3dl0szgsXUwNTNslljeVoImU8
XBTdWh52tdXdIrdtY1WL6DF01yX7jLEe3ZuaY1jDzDkQS9uuEsPNorR+udH00az5xmvyCWSp2MMX
EnjbC7emQ3jhAMgooMzM8aqjfCsTPTvFTAh9TIos/ktRhN2723R4rKr+YecVVAr7nBEIH0FwWA6a
Aq6h5qkQ5cN47XS8dsVfp8renE0DI4uf9QP9x5rVMzDdd1MuLprQb4eBbQxYxaV/8LKctNkCAHTz
WUHEla0/Zycw/Lr1o4Wq4RLxhIdEv6FBWqfe8vflL0mg5iZ3sUCwlRklnwPBmwj2CnBsjnI1pKsn
7JHZHucy2zNv/V0Mw8aq9YvoBgS+cPIAkCYYBFOY/FJXuRy/R6woQM8UJV/niVXZ737F74eXAYJ4
srQZ0QwllFqB9XprW3+ljVJK6E4TU440yN2BjleeLfuw43qvlz3Oumw9ZTCLkdyqenqCPTYAE/7y
fOp7ZsvabvAVJKPI7bWgGJEdqLL+Pi5lyRPFQu5wIpoDaRKF1qk3pnenqAtrzeo5UJcmGyOfcCW1
BRgtwiSrfoiXy6fjXAW9Q4TXIoxmlAPE5/xflCLOpU+roYiSp0IfD7viQqZBuaqbkLcT25vyAkMA
SkHWBNqkoFd1NyDn5XIfcbJg/ORl7ARBpSR1zO9dHToDNzzGhZNGsgjb+az16UAZ6PnhomcCa7L1
84QHkXFSSzp/A9xorNzmuHChvfUdatG941/cWeks40rZfc0kN0Bx3Xm3HWWwyL+FbZMshkpSGCJ1
MxzAKNofaAwJ1JuUbngaQXhoSzMl80fDiRp3j+QUaWxCmfVed4wh5yzhDxMJBG7ABspH+ylBsKBi
yDRfI3jgTALDrySOm6/nX48I7TcWrh+vYz3RPTHapBsh/WVqcm1EmQ9B3Rqn1mx26h8mDsEAi/ea
KG/C14feCEhUOikeZNBnJX+BZfjl3S8TIVQwHP+NB7QuZdruaoDNr6z/WqUmzVmNv843/DPtqPYB
7W9x32G+pr/oZZKGt0OgNa8jMUS3xgrXrT1gAw1zldtIDGvCTgCvS3PJgi4K89CugKWPMoE2IuJd
zz5P2aUS4yTv/y0gAPRBUcetUzcwgjzOTlhGZf12jbBoG5ffF3Bhv/cWo6/p+38R5/BYRFu+ifKh
UaJPAqLa5wSbTIgKnFAlkyx3BV8vzqCr6zhJnT3IQWlhtp/JS9bcAfXx+o+6y284rQonWqlRItVu
wfAstQiChkqNWuLw3Dml4Td/TNkomBj1qdlqpQTe2D5w2lLqPdmagCNTJ1AV4coxsVVK1h+gg5P+
oFNMP5VYNcDm5TKtPcRzR0JoqslXNtCd5lC+4rIIlZvA/uvkLydhzWkwclAUZ4V3dngTsUyFsXDG
f18Jv239wqrwRtkDGgHT3M3s7aGN7is7f7uTcD8Vr0GNCJQTfJvygWV06fP+RPHOiYn7bFI6Ov18
C3Cc9rsFqpR7PeQKmUtXbgmAB5zyKxN67oa4Imk6C/pUBtjOMZcdIEv1OIQgZx0uq42T4vNjERuD
0fBVlREJzIKuqw0/hp1aeMRjT+sxVCZE8Gw6/Xan/4u9vnX84Y+AES2fGt3b1Wk9SeIksckZnd22
qDPJa0di2IQlWJTk7TlHOs7p1buGiktN99ritUD8xPoiBYEPZ0LbZUqXHxdAkILjgwoByWut5TZ+
3npSa8e4uOst/nHxGmVVeZtkrZoXyXQbV+Jtht0qPaD4sp991b0vFxBsTkUTUkPB9wd/V38JZFPy
C680qm6awLBNv4i60cvY/32WVHT+cX99gTZT3lp7uzAreqkh1z/ztKzBonoebodzJKXFiSovg4G/
DGJ7rONmncC6ri8y1ywe5pMts/SkmanysqAl6uOsnH8c7ExLQRx7hdBFpQaTxbcbJ5Ss8KSt6Rji
NL0hYAFNZCzoieMqhcxiIKrW7RL8WDT2DBgY3XAPpwBfX8UVIHqb7hdvWW5oe59FJmxExnAjc+E0
GbpgZS8AoRiFrP8Jp5SqupFj6iFj+si6MkL5vM1CsOHTMJXn8DJP54q+GfiTfYz0zHrTF3bWR3qm
m1SFTy2pU1v51QHipTdiJtOVvH2k2QcbKw2qJhmFHALgmVXe7tKi8cLjRU3BQffd7U5Wx2ez7sBn
p3DU5HIJU1KyxgItaBMnLaIGdvjArFdaDXZYTux7mdIH8fd2b8XUIMWg/R168nDQBvXpi8VW+OR7
P5hcAupPC2s/F7qKkAC63XkUoJlL9RaXbryWp0RTKM62gl+I1sJPxWOW0ygPxDHwEEbR+7bLgErE
hx5BH+fD67PulKNnpuOR6IzaZD4f0Knz3NsDJM/R2tqxnCyEB3LnidPi8b2/vDvkQEVD/fUE0ore
OkXWzvbWjru4/DjZZxikcio3VciCOkn3WU7BOZ12aciKkUsKUC/RNgEyFDCjhK8T/1SUey0RpZi7
7xVjtznxw9Emakz10o4EBOSXrrvV/6onBktFQd92hdfqm9fwn0Zl1Gx1RhsWy7++dNThEgvt/xLn
S3JgNTQx/jE1PoBVTlmWqZ9RbuDpu7OsxynAqUI//VRVOsg6QZcK3SHNtrBZfCVfwz5/2KLMVTTS
k4Jd2QXZA/mWl+op4SyT4ZUdfoMUq9QlTGS42KSVEajkIhC/iP00I7uxo8BgKh6c1BXAKafNEjcC
006+uj2qn/0KQoYdpasSXU5PZp2P7gYsmcPPdPAztMfOOJX8QH/outjV/ImvoakWrM8KAo7rxvdV
LYkV6CWjqTupAI+HOHRJdOog3ixHfiGMcUTANOtdtHnS3nTTmbndtaqIDQW/qqwTejiv33mqalrs
h0cDPkW7n+mKjODL8lwLxoe4MnkcCcLDsYjBcg+IECeIuSLfc6oy1J4XCGLxHYd5wpWoNnsbvOHZ
FZiQ8aqpOHboyg489ymiR+62N7X70P2A7M7Fax0DQyl/KXFGcqvP3kfBbBdtyVXXirmMwynyaZRT
dPrFQsMjA32ztMYzhKvgOkO1juYp5AbYtKn248RddrqtWgF1OMnoh0a98elGBrPvloRo69WPXEid
VEMCOi41BOh4SDqyEgfauryCoThdLksYhcQJ/F2OtHkKayGLyLs334CHbFCKYKjT1MSwS4B0hg5F
qtCWc+0S4gD/XAOZ6X1aK8muIYJHEwkK+Yw0ADRlipvuHqxM8b+5MwJdXcdx/v6wBod0+PvcnDJ5
84UP71g+cGP/1Lg2EGzlR+iGXihF7QIXbG1v7jtafADsHJA6Ktw7o2WgXbad7SOZCIYTXfceCTMx
75T+CpHva+ngwMjxa5AxCC/DRMmlBK/uty0msIlI5sv03SmTaRbZGCYEc63SFEfn+ToRsdulPQvA
idJ5WGvN7UCzyKeMo/VPWmHCgE6v9pGp3lit1TtTTmAUnP9/r4APcRdrTQVhukknD1WceP8xGGT9
2Ir1Ak4HiX6k0xTLMtCEEuCeSH2OiZ5mvyI673L28nkSuhuyBdacyxSL6KtH4Oj6MtFQmCWHO5jQ
KQR9WwhqlnPhOeWut/y14COzoGYt6AKAD2bY1dwck1RoSQDfnk7wkD0RKenm1Q0DGhvMJ1APwmmp
qJW3tVtzgdXBA/C5ZA4dSDeAp27o/051Ao0o/ABFZyK24oNQPuvjeS0PncdHkNevv2zccolPm4yG
4Dkax05v8wxVSBa3xsDOZLsJL5CZY5k+3HvMg9solxEm9GCMgvk4UGQ1LuVc/5eFVjtLvexGamUn
PxXNQ2qBR74R3pksvOyP61IW1nwYC7NzkmwZeG2E3Bv49px3JMNjw6MEaUBNeDQtsixeTjzHRgyz
5KCXTkY8JW7vs1dU7b2pqButqw8wOwLpjkb90K52UnelCQ5Aki/loAN/1kN2lsp9WuDcjvW7Y9ab
zwusnsx9kqaaMDUZg+daAGKxp8Go8RQTMKf/9z/0Q5PIpPmBpOqpp7f1yBKLIFbmlmrU4ddExKMx
nZCNZ+kzQ4zljJiHPY8/jMcwoDBzpkU/HyAtKu6dGslVuc1Dm3hq87TQ9/zz5IZHJNT47Ld7aAKr
TLcPuKAtS3lQcvQsR/pyHqMnFqf+8SPr67YAaVxls2cwcq0jN4xh3T28e+TGxJoWB0RmQ6TVYBHV
nz67cZxeNP1et7HSiWjPEcPSHet4kuNpPto3Yxw2of0ANtOoExPYqaddYzOM7sMglWQV23ggS2yR
nWheMVURRvIAq3ZjMZKITMUQYX9bF5NKeQ37BUHMPDVhbco/3gn6T9mI3n6GIQg670NTjARAEmNA
QOw0yUGbhujMUd56bdDq8tgZ51CE/oKpytlJVQaUkwoDIzKiYkArHHdOBvKZVQfmDOO4S0jQXt/i
ESjK3yyt/DvCoiSUOmh290MyA5nS6j2oNPYk8bOudlKnz7C6ZNMtcYTfdwiczpnGgbdpaGVwtntn
1fKnn8jey3sOrbKBfEpCnl7VFpkn4QZYE1chwYGr1R5rW4H4/thIKhWKJA0StxT0UQDyBmY7HVe2
IE4JdAdRYNfdLJVoEPaNi3xTZPTEX6U7hvskTsAdTjdqV7aIet7LraL/kfWHtMFseVri7lX+powo
d1AbwMXyKFP1RrQUehX75PvzeJPWK18A1LNBC/SO5ntxl33XLHwQa1Q+yo7/2UOGZ5ZneXOnFJfS
syR14dAUj0+rm4p68GDnmkiML1Pz508sWU6nxokTZP92ekpcZmXt7dsKNl/+B4G8CmLopheKHfZZ
EqQ93sVxILaFTaqy+0bWOdelfVMrbbsuFObkUZwPiMTgvuFdKGFrz0yz+uTILt2qqD4N8sqZolbL
kxODY4LtvHfdfByLDUTkTKkmXOVpF2FLM603nznsOs+Mm7ADhr5FncBbS0ZPWxATyESnHRbsBzM7
0WDWiJ7FMzSvWdI6T1o+xm5IFOGahgWIMutylkNzTSmCe8Za0cKV7glKJCtWsZoiKnFwHLl8n5CN
uHJ0BTqOEgTx2xyG44qnDVBOO89cHiksDL+7l6/BxOt6Mv5ixrMXtZaIVYd3MpUNWZ5K4LsWJszl
H+0KfmG9Tvz4w2+4YhBycDFhOalgaO5Y64HQfK9JageVh1E13949sLyN54x94Nv0JzBeAjOtJCCP
RQALFbcUdaXKOqhiLrFfyYg+09z5vqDTPxuv2hCOZp7KrhlFqa3CSP5zwpMo5mwirWC3R5zSeUC4
Xi/9mlh10JYnXar5LfXIc4Kr0R6OkwFUJd4fLQc3Ns+2GOZ1Lcztb2iiXyEWhc/KB9DEYxTAWSB9
HO9nrZPJoSFgR9msqQCIwEL1287P26JoEZrCydCRyf1brMf0hpNtn5tiHkGUTYdKt+n2X0id3i+l
D9npLYCnlOvHyeNxlkEi6fxI0Qnn9kLjh9r8LyRKaw+jM1lJIupgwEAqdLHpvIbMQbMqzSftqA4D
OJSVmdV802yZNuL8S9eubVhyBj0LletjME5E3b+knTGXZdUO25qTbCbr7ZQ+xYKi6eDp6A8um27C
gpYrdjqU3ng/y/QQF1Ml0K/qfBCQTEDL04i31g6+grl09sOh7yDGrLdvtkwcdD0ZCJNrbxFLBatp
A/xKmQ5TTF4ejv73kElbCQa8VKgfYS56QKCeRE2hHQ0pgeTDHcweju/s3uC2JYLTzZebmgJKpk/B
iiU4XN/FDWY3Xh6bYK8Z6PSiqRaWv1WPkTptodjUZHRbcALiD/UQsKIIJQaLTsXZ9y2kWW1CAZzT
z6prmS1SxiW7X0R5+DmiIrclsy7QfqaRL6/L+LBOZSwxT4jNE67TTX77JZeu+lmR0cbvzr+0GU5K
XYfuYP68fGGHLN83rQfemin7jHoiKhx7/4lmTrMSzrWZulkNJg5VSsj0QlPYKkia0MeG0tod/SGi
Pi9Zp8mUQGfJVoyYqM6dKJFIRr2JntP9PunEqHIsF+gWgegzhrOahL+PUKs+Jju7zqsvcvNSEJZ+
PqrU5VafjmM17iQkRqNoEPFofToRtgL9pprkJ4xofqr+2BidtMy41mlloycjK4nl4u06VXqw8RHC
S8pWv3jcf/KDSuaRv/YweFq2Fl9yAxOzGZ/0hmGA7ub4inELEdNsSBvG+LAxhu5Jl4TbqsbVIFK4
drZjOnkpevuTncKdeg8RSeqwcDtbaBHXpPWTX8zodFpK85jwmVULo+ckMFMoJKtOspuhKRZtD0rE
FxTjEF2L49DO1Nrr8o/O4uBO2Zivvf9Z8NFukCOfIBQVI1I/Qz9aoneMDwzmFAU2TRG1l2zycicD
OLNkFrdADu7cGySaG/EIhZ843cNdk9M94/wRk0J10bhUtpmphH/Qi3WLPEhmog7GfCpfclf0cb03
37qjIh1jdhyjgTsWJ9oOtMucPG4rlH4PdiVya037La94WtyfMZE07OipnePSagxxKvMCD9M6bnNE
CtoQNkrXDafdpgyxUr2IpBGo3OugOaGfCJWmZmwK+FL0Mk68atirqEsD3w5tRk5W3qxVtp0ByW6m
vpSvdnVDxpERjndU1x8exF3j3nB8X0BBSPol0Xt/geCDkjcZWU2E1cS0y3V3zwbAo0+/56s+8mrQ
Ora5yiT3K0SxQ1HE2wims/fX4rna98hFZ2za8FjviEpuq6QwBtCqAcrbKMZuIyo3Z8bTCU68RCrM
VuVtrGcHTxvLhSBnLXXquRSgZp1Lysqc9pn0B6oJAiUluIbN7EjrMfY4IKegFGTyayrObzQuvfqY
WPPfRFkazEEBpmU5ZiO30ISCh2O8gQ3u0ppCEiWLVDFWYYJW3s9VY4cqEsBpNrL9c+SjpzcmowEv
SS3coZaJJtjy4RHgQyt3gQuN76/ufOnGag7q+Wxev+xjuUrjwOMrcDRqlaEmeiPAHSR1ILJELINM
KIBJJs5xxiOdGK16MMtnihN6Qw/XyiZmb00QIOMZ7koEouYDtGTnXFWCgw87JKZEkTJfyYBW6xHU
JArKdi8WItUA/jvz7gs5OhgGmausmq4UInbgYvYCXQ3A+ahkFHU+QQQNVy+JJP3L0d1G2eojL8QO
AAQ+lk3nPRarW0SIp2NH1vSeKL84etwbrkyHiklI5Hhg0jQuPmWvgEt613VinY9B7IYZSbevfsGU
4OB+k5x8ZGj3SuUrXPmPuxFt6hNtY/DJODq4sMgCaHTQZWIt4w6dn1tkzwdq5Rjp63BHlzX47w2Z
APBaFdnzYqSit8FNANtdPpSgWPEFL+3puVRazPnwJP1mQMdoYE00oDzZdYVtTKvK6nGQPxC6835H
dO3/6Ey5b7mZmcwmMRPjk0YVc1pklIHPG2kaDtiwAfnf4o3HTDSg4fOK8f2Pc8oSBLsKRnbR/6sB
uMKGP9BKxADWZjl7rEJbcjdFrDXVSTXDnnR87SdIYTUyYLJA5Eeca4IDUvuj+ciOhY1l5XdB/Pkp
inN9TtUh0A4iX+alsf5JulI/bMBwQGSQeO96M22ze+LflEk4rA1X4OZRmKjOynYpc16J+NAss57+
dgkwb9C/p3JTJXnnL6FnMZjEoGw6qo3SsQwI5exSWMYhn6UWmPgsRDYkbfK1lE8krYR7rqvkJt9S
8B0fS3I6nJJxNscZU6tAF859gzcHlCyPXbB1CrFCQOzSceWk8xNFmALLat79SpCNJpE0HP6BU1ju
uEoSCQQYlhnLsHnQhyimvYN9A28FbieI/Zy1J3IV97uSnXF0om+/dzdNlA4LNyYPNfkxUi66PrVB
VRfUl8ijxN/QMcguW+W8qCbKX8hsnqzF5sPYNILgpe6HeG7Tefwh8D4wecTcC+XCMv+wP60SjQO5
s5R28CLOegTx+XgPA3cw3gW3frNpX1mCJotR7qab5MiYkoca1aJdLziT4Xw72oZOINPtzMABSISW
hLCLvmqz4Xa6BPmJUBK7dc7gNnwCA+UHSJJV/EbzCNafP0tf31GES3h837Oygy1smUtTNQkbVA1R
t+3uvkylwOeKzHxf9v+7ci5E8lko9INj2wuEC3zJsD0NS6WjTZNjgD/CfAORiSSnGj+mAG3a3FnD
DbWVzhkoZVRlduClppesBcJguKGq1paK5IK8RJ677Os9NCTtemCOedczsFYazl9x0CW8m+7wlgGs
jTz35scuehD9Lt0erNwROmqwnlUjlDfe06XMhY+uIiGbVwvSdZ2QLy4x8vzx/1TNFs/tHF1pEnET
Q2v/AG6yo3jA0ILrMQnO3vUsWUN1rKhFbZ/oZL0eegx28sC8kD4qwVJyMORlGBLj5Z12LVZtff0M
R54vS8oRa1nP8oXx45nvvAYPfrDt4VrCNUGNkAoPkZKSKkl4jocbHMShpAfdz5dwmA/WW44evVcj
VilVCBZ+Pevw7RmRFYPfIEVZ+IfTm2HPgkCXTSrFiO8IAHqZEG/8OC/JfI4iCJbtz/WqscKWoSyY
G4tsPMLYKuH9yu52UVCCE+M7e+W/2XAZr/0EQGOEmInuXC1EluLaVzn+FHHjFtVA4vqAzke8ydDg
4zxcUF8GEwBNJOyaxntAjrlFDB96Ue4uUhnb8kVbd+STzSf6hJcKeJVv6Ugz+XAAgqJHRNN6M6Tf
fCFRhMZJziRtZauhNKEE1bknIdZBpRT/PA1c2M2qiD2IG7kho0PUm+/uRpHjiqaMucA3zE5kCxNP
p4KsD98sC2vkPFebBJCbcjw1VUa4yMBPa1M+OSRgmBcSEbR0RBFKE8wy1EB9cSVmL7/J9CbnJ3GV
Ye1qcVO/dnAAqXJhji4rnH9Md5uWWtuk6vU+KGVgFxkSc7DHqg7BIGc9N+2p6/9xQy0nXZve3doe
9AQ1y4LVg7ZoiP9hfpqK33v4wtWZ2Hi0a8pWI/tLokZJMyUE9D178q2byqi8XmA8SbWO5qnkEyNA
JnuAO13XuGvbyT1bwvn+9R/UGOq0yIjK7wEIufIsc/lcpEhHXSFl8FREpOL2Bc/bTLJFdnvzh1/K
ex0/KCI4o0fal07hKmP6v7Kmuy89f0J83FM+0X1bGE7SKOK5QwdbL/h6Cssye6KL8X1HIncBVp+x
icFXnCtnmkExW6EF5ztnf+97iprTGGl/O+kaN9psovtT3BUVt7p9UeDmB2XJAb/i3OLYHSw+SAhY
74i0swHMaZty/GRp6LC/IRc5U6gM6PP+qDCulI21s2RqkxcwLc8e2G9xr1p22f1wOn4P+wMjkKFb
gZDFGikyqKyv6z1yNsR/fDOUCenwmotAB/rJF6MzujIpi3YGhcWqgXIVthm4uUMFgGw/pVt+VErZ
7DemlbPz+eKD3XePSoelPLO9CsbPP8o4JI35iRkcKPkBrdFsQgXPcCuyh3q1MeI2DAWKBfT+UqSK
j6FtIzvEWviFQuAQBS4ynMUcry66HmsaFXye7E2ngC3p1d+Nx8isTO6uXt/WrFXQePNJsY8Y30Gk
UPWnje7nvM0YQzXDB0cTT34+WQWtImbq2/HbA6aeP9/hBAemoHsSpt3YibW7/IxiLv3Cd9bfCTVn
F/kyAwiAI7dbb2EnqMc0al97ZxDy8d02l59ze3qobKTAhQh4bUa/bTwuNBiOQAO7tcPN031WUGMJ
B9SFU5QEakIQN9Gv/nmFliLYc0Tfvda8DGBpNq4Dv+VeG/dQqu6cLMiFSkN9ZpYEWepD4b6WOESU
YYBH95fd1P/88ch+D1Sx4j5LFGAQmuGvJpU1Ve9hBGww8VNVQ+gi+29xNME+rm3KXtjr5q16+QQv
OZ6rTmPIc3RIqelIUbYsOpflfBhB9GmmvlVcFpfJswA9SgvZYR4AGv/atKUA+B40h+bEBQ/9v01V
N0lujcYVCtEsz7SCbTLwz3QQ1Leh1+xCa921fwvueEy2Pih70hExIXBC45ITVzASKsv9G2quE1aU
oPreWyLFqnlHD5shnRjMnNeUQHE5yC6B7P5pyCDVDBz5QQkNSUV8ICmQVJSNvMfEyuDLoHdzyTn6
Pmkp1ETFn8NGpeHOET53/3BKliom7s8lT/U8NLINZX7R8SiBH8mWmfA6ZV4iaQP+ftk4VwStcGp9
w2tQqdQ3/yIf5iag2cd61Jv36/8Ad9x9Erk1p05TXdMeCHPzvDIiKRD7xiqDBKGyQ50BEiNop8uF
uf+7sYQqUQX2COSdXbMay2XjD94AtxFMzC7H/XNUWyBCUtssasOacu35F23L8LkzvHvdM9JaJ4tO
eyXJK95nIq5t9zKSbgaCqmp6GmvnvhQGGrqRhvtI4wqZml7bSZ23RIPD1n3FKSoE/xuS4Ck00aY+
C0Y12ob1g2krW4RnyrAPDlBZ88fCZTJDmK1kS59GJhsYp57dIimSOHhB4VSbqAm5FVpi3RYrTb6b
xptQzvuJEfBpAQv5ZVueojcfCwLI8ZSBOKu21QRMR3A3klUVpfbpDEHLz7F1s82pRSngXmjF5MIW
XIgSqGkvVdgMbEsyQHkZEPXdWwWaC7mjtWIrNayf79pfZJ+2QTitpHg0gccY5F1gjcs8+fXnLE+u
ERzfk6Ndf+KbF6JYw1AMDUH1hCvd3YO2ftatLSx7RoaDe2TOcOqWNeXc9siE3DZqYE3tBgEkPY5A
nDB/wSlT6f2ShiGIqjDD+CUXvwvraN7v2QzUHQcEMXFIdOmj8p8dFwU6uI3Sok6ujEwwgVsV8Tzp
U8ednHskGZzvOa2lgWtD9nF/CNrXNhVh8GzKSnr1pHnczqr4gGD3hL8KEWsJ7yqPoggBRw3j2bW8
HXB+9h6F1uPRpyKcP5m6xPEETYNpmHQ8K9L4xIC4dRm8IhC2+vKyZdEPghz3cfrjmGU3dW5DXRi1
HcsncS6xsbzsWpja5kSVjVwSavN5ZbLkReHBqivFj/q2issLLecb7T+Y2MI1sMguy+T5KK8rpCq5
l1sbk0cmJn+0TvhlPgF+CjKk9a3LQ0vuiFJtRhca3ZzJc56CQ12XaLF7G6NZUWolQPOTM5oDYopN
LJ6PzwgV6iHrcu40OOpW06u4xsmWSFiyeIRcPVhrsDuSRzWDup4rT4Wg/b6/TTqqDZpRvU8pUJuk
4Y0cfk9BKdUMAb3uJaIOUharyx4pnGvCuQ2I1W6W13Flf1GIngL8uuI3HiOr2IRiozo/wedB4rYl
sbZeUVzBcyLG+j6TFwkMJX4LO4shSJqKSxkVciu1DjfxY17dP2UJJHtHvqichfX4MlSax7vHJz8E
IRDbLYGI/AMU+U7UJo1Y9sJvSECSiKya2rr2QRfkUR68w4CA9pgcUNZqproqtOVG774uZSCuEnSb
m8CPUK9YWDwfgNMzaFenImjpLjTH87y9inw/EmVoN6Sp38lJMK7C4RnTXXPzgPF8mV2kMWeNwOLw
eIUWnayjYPX8LfZZkWqWaEVsceyLS554TrIOGxZr1myefbhAvCG+/SDrb5sYCE61uMk232DRfWZl
r0nWuxy1gVcMOPq49fxiWPeM24+GW2Tt7IUveDDbY+5hgR+47JaTYdA/Bxlrf7xBtIxNHdeE401H
4bTmHSOVbBAZsfwP3vIMSceIF/ReNXPq5LxpDZotJyhjgr1tq3G6Z4EmTjmHvkOWBcDb7ujrgn53
QLGUOJtf4CVRKpXqYHzYcTDfYrRjXXXQlv//W//GEsO+c9fwOqYhqmNne4feYJSgUId+uVDX5VKH
6CRh4EMfKnLqJJTnHFDslZjfkgyzxa8+3rjxl3x7t+wRpWTpa35h3zK2JQxHfCuoPJCpHfjoHdoW
Izir1/f1Bikw98FS+Y9WBtz+eauM1EJVzGI5Q32GQYOrTRNjYPC33+QF5U8sD28P440JubPD47ba
li7SCjeODB/8ZTNSWdOgH4t8RIXDbFfvenZ5BlJ+2VNUWcqWE/VEv7UZ6Uu85DJgmNq+b+nNC508
ttPSKSx0VOQUgLJoW2+DDEeFF0phWaCopBLQ0FtYS3H/N5N0ynerrgaHZrd9AXeUW7LOCmLADehw
y0a3TNMA457xLqPMJcnoWwK9oNZf9hgL2Zo5b7xYh/6eL+218VxBBGFjgWmnDJQK9++WtKPO++Gy
VZrD7PvLPD+U/OBOqb8zyI/o2m+gG6TmZIOlkpWCfcXIBPftaA3EQJtJq+c9AgFyq3789VmfeYn7
MCyWgMQdDgcG1voW+gmaaaan8CGr7WhuOdIQebd9G8wyBaAvewZVIhjlw57sO+mwfiXDZlIXrw+9
pH643IQrPVO7VrRAZpp1TkcXRJtL799DeXPVzLeLDSW50bir8voNRnr2cskimuwxUz7FtosncR/l
lb/36cvc5SMKVtiAArb8TrrgLsytsCLRn/gjyv5BDCttZP36GPPv5Q+qrh+gvbp3qaCvhs9LKsJ4
AuDAjD/6EfsOx2671Umcyrt/XcKagnNNf7V8zOaZ1GO4oH4l6gWLfv6Typv9UnkngPE5ghLUP1dN
jLiECmcQO90g+XCeNx/rcwCt0L5XtGGLpyOTWuDneUA6J6zKA9L4YnwA8uR5pHT7kJmmCMDGL0PE
98tJTd4Lf5JGIpNo0rA9zsNCM72fwwCxsdymPk2r/8ZyUnv0SeKYhRUzC7dKnTiSVoy0Y+l9aA/0
xMQZOtS1tbcs/eWpgfQTwZ3VsjTVI9j80qp8JzqtJ30uJESPQkjsHEYYJhX7ThdghQpxdpl9r/+H
s5FH6Mm+oCUdEaOPhV8svtR6mjmSmDxttLTOQbyT6G2wlDBJT2Ax0M8p4qZfRNBvofoBb0L1TRVl
mnYzy6hQie7Ddx9D+cpVVJpdqmx6a7uVHUzmX/1Pc0A1wFXPNGphTDQ/MycRjsOfgdevJUfMkK+q
x113ODWu44bqc50nuTOXKP/baFfrhrXULQwQlvbt3E9JRpWgPcFK4NNHxxQ6b4EJHT4ePG5txRm3
uRoOA1bLh6Th1dXoZQnRWSK+2v2XYFa0YFKPpdCWIB738HwekeFjipRYaLsTjcD5sfvIfMaPwW+y
eajxrn6bxn/GNsJCXEhodQtrgz/ZXAA7RFyEdnv1JPWj94jgV6LSh179ak4kym1Ezgyf9Lvx9dPi
QeJ+hIf0iT4knq3PeUhL20pq0XUns5kh4LWXWtaBYOjwO3GhX2Dk9NyCaf/l23qdVXMNt206U7AT
kOX0Bhk99p18HM8BVZ4lz1Ck/Qs+LNzMxUsQNWrwHZcj24XQJJbQXxkIT9gxPLYGDBfsu8D9oJak
2+fzd4tph5A0Db7AGq1reJ5mNfnI8E7KoxHQ1CjaHdKsEpwIW+/18yBB9kyhIkBjWUGn/d6/zevp
neGKUTe6l0hRyQx0HbTWOWybxplPjb4ACUE8FDPq0lBaOGVzNVe61tvuVCh7EzYgQwYTaTxTaXmx
wii/ZHY2O/2KzPEyuqyQWOLtVk51IbU4OWwkaDlxhjbiZQhoEj5w3vgHSKw0VyCHMrP2f2hp0e9A
tjBzKJbuIUMl4N/3irfo/CbC5SkGgB5EWqgQ7JTpShmQsgsGUXNJHp1LxHNedtEZ3VDxG96OCH7v
j40zj+8PBMaSuOp+tjNsIYrXfjyzYc6WBlCqSe2A0kLPDuxmCghPc/xqyWgNmMytkjDHoLOZVcuh
CXenSHYkDu0SqbDXbbiSwtSJ/ElxFSjHCXKjiSdB05OpnXwUA2N10PszH+bXRN235YGo66LXM2K2
CRDdLCnD5ysPGHCwUrhuVZ/1xlIYu7X+gqdG3uU5EfbwHluahQRxuiVfAcmIPpNUeHW+MbsigrsR
IY+3APSHrXAdPvlJxyq3//ve4gf0WAYZd5UWlHhrH3yI++fnqIGt6PK/stOh735MrsOk4sEwEs/I
AC0xDW+84V1XzH4XeLR7MXQ+0NlZ1pBY4isqV+z8jS4sXZpIsOpuw0Fx2KAKDvb7JavEfUxb8zxt
oE0xRSMVcTbvnyJn2DS/+oCkFIxDQ16vanWhTqSuY5qgu3PNR/Rydu9MnhPGg9FqDYuKGJS2utrQ
1c2xzJTMjGQ/sg4EpgE6kS0TJswsJ0GKxrL9ni9M03g/+HnQRoWTYVkn92BwTM63NcFrBwflGTtW
ChYl+PnQmdgjYkg99qP4g5+gZeecCCGElql14gy47NwvKQLo5Vb8qYqSvuFOw+x1xu0V5vtYZxAl
Y/+BSTLnxQzNnsuN0liqJ3LCwCQUinrfNTJ8sEPeVeNXZ8xu9379cjEzwtKj/bOn1jWEUxb8Q/oi
2vBlpQ9N0KUTdbKJZ68I2Gw6oiTB0xtYk5y+rs4PuvBHUlhUAt7+0mtB/hxrAtZj0EYXql/e240B
htlKq4JH7vORrLhc72n8KmrZZvowJdwHwbiZkFt9BjjPDxdD8ojtX/SdWSj9pVstNYfoWuEJsPlO
kbiuDFebUvQTLS5FXO8WKAbg2i9jqH2s/KR4Cc7BYk5iJ6aHubjd3kV472RGgRWN2JgjyJOR6GiW
EIWP7idHUjvUj8yTQ4al2MSePfaudz89d5WvTjRCUFoZ3e/rTYnbro0t6EAvGvXOYeZj37UUQc2b
cm4/Oq2lksXVk03BljZIAODLlGGthFlJaeyhiBi6xmgHuByHesWWVK/0ifWMk4O4NltvoYXlhPc7
FiLfSA20UVO4kD4k8TFCGFzZn5QchSoEogx1vsF6Nb6xHntJX0uTgl8K8Fn8FIweYIAw4tD1Myev
aZln84XE1FClNoBS8amzdXDDy6F2Z/KuTHtNzQPsIQfU1k4NuKIP56LJ8KJvlThPc4WCykE0ZLr9
Hq+IDGKbYc2UseOfD3oME+s886KQIfFgLMhZXAQz7YPGlW/hLYJ3GTTMGZWtL9DHMy9tl2dtfW4b
0O2WnpZiHzd+ZjEyC6lOSIliv0y0cNm1GbxAfAVfl+mSZR7IvuHTRHkizYlygc/+TWEsnmpNU3u7
0+p8xFOKi8C8Xche+lOdE8XbnaqA0Qd4dzRo5wjG7/hYpIVOoV2HDq/m0/9Nlh79kdgHyNOes/HA
Fk88z8339XtbbkdjLEo5M9PSZdNq4bCFrz08ZaNFGDLIwuMXDuIqo5/PHmvPBj4ZfkcZ+sxESlm0
SThWumvHqgurJZ7qDaIGDnVl8l0KJfmaRAEQ8Y5jpu5v6cnwn/BctRSn2ioeuKACg6GE5FxONgRF
UjLLXae3kZrcCwl9zH0ivV4dlLYbcxd2l7DSzCH8lHOD0vole5lTp3ESRUAG7M/tBr6fhgzi/wFl
MVddhL40Oni0P++t4iPzrrFh81gnk55g93nQsITEMT4GrDPJi3pppUFSJSAXQ588g+J0M87AYZVx
ugbMtn/YEMyDJd1ztneaWc/rqXIdessfuqfNaDjL3Nn0ORrnuMTtcW8YTepr8QreeZsaLfgxRSC2
X3/iTavyZXN86eNAqeRQd63/Mzl6KiHzW9NgtR3cWi22gqbX1eU1r4QFr9LepooIRnt/qEmR6PQM
wzkxt/KwkQt8GlmlbE+un2M7vGP+eaC/VHvb7+Av18E/4w0TaubsNpz1F/Kgd6NAzNTLSMFmsUOH
DarFLEV9dsp4JS0a4A5+yEnGlFZaYRDe5Dg30h5L9MgRV4FHxs9y1SWm6RxW7tByazn1NFmUG9J/
0LmgiIstWR8CUGaVOxhS+15K1mr2oMSZT6egV7mGghAWqX9bM0QtNlROFAdYJWMqk6TQKo0wG636
LUhSoBWpmLFFDFpA+Jpw8A0D2ashGmUP6FUkeVKnCsVQqtaUAVYXqNpbbRhhCy5J3AnlaNTV5JBF
jI8SBx0rHq6j2PZA3tOi0AthihBP3mU1YatkeXmcyPpQFedfj/xgLB5UaqPonTwfTbEhEK9ptT2h
dnmlzdiQJH85l1ASUH9ov60hWXR8PXVxd5vQnIZBOoQKnuMJv3qvvYgk+FHUxUfC2EHBOg9IhmZj
WNG4FuL4ghcGMxUCq383/Zkr5oW+AKPnpCuwyecYuqE7sta8LXEGK0LV7bjW+dqyVdVEbyHLBQ6y
D9/2xIRp5sNi99n3SZEFVB1KWmBye1ngvD1coVR2pBEklO2/ukoSkpW+TyGMpJgFQZZnt476h1wo
1FpwKuN/8c/bXAi3/MREyMVrSscli04ga2BT18aBqJWanyXB7L6DmOyGZ8Dm3TqQMNsKWL0GE6c7
JI2QDI1uLSdyGBcOvh7jEotwWw0RZt50140cnCExvo/0+vj9PFxmqVE53Z3b27dmOiepY9hUeVRi
Gm9fVA0WiQ8ofREy5ikKYH6eyzTVWKDcb12WCTZP84vz0tUA8qDIorXonq1In/UQXW6e+DxFiCG4
57e9/SodedTufTmYk412lmMJE2/6amdvlgbcACgbVXRZ5iD3jxThf3xJuLyhMM/1dpzIjltmDhXq
a9ZYQftPhbNNOn13A3/LO0lAbmp35DBf1gHUNP7Ej88DcwFHxhO8TJt3gEVFLru4gGPlnkD4cgva
jJAsoLr2EttLnAdEADHnyBYcYmgTJh78gVzOivd2/KA+3OS9R2gCph9n33XoEuB7Ol/IpQY0duSx
mfeZpz1DR68cIXDeF3w6p70+GM6xArYXSyGO/CGiBYdSVa4XySr3+R/QZBZugpVA0smz2lQQ45N+
ySv4SKaURaZKKZH9HtlTrfz1RpvpDI+XIZlR/H5Uioe/o/0tleLTClIhpGLwok4kIrB34OHoG23X
tffZCeQB9IMoQa4M6l9GabsKwfIOhP3Y2cB6U+dHNC8eF3PlGCM3ZLRW8O1GRqAQUbur2VM0vegQ
G15xlTENN/R75sAzOaFLx4oSVb6YZUlk+07e4F5J+pdCYSluQu1DB3K1TQYWd0MU/vV/5r8qmM28
VNWcOW7eNTB/Lq0Witu+dhIgwpFChGdAotlBgu7gPLa2oowfYzeC4OlKyuWPlmyl5QwH226FVGsq
YRM87QdrWVXS9uhF+gWCpFZM0yh7qiiQ/0tWB9sPCqwOiKUY2pQ0YIhJ7lXhA9BIYqT+Xz2o9yn7
G4Y5vWHVmxeMEQdq1Cqvh7r+U/l8ht67CCk8WgUpL8rqQaa6vNSJaojrZBnYyk/VwJf8hoDoDG5N
h25OJFNELVO479vEeNA0QF+RckWWdODWskgHQYpVIYygGPsbYOr1a55FcEUjyFLFJHDcNADF+FGh
hxb5r1DrEQe2utFriYsRd8Zaz5dIqtCHGapG6LHJNj1ZESX75rijMlrfNHu/sXDrJzyz4BzyJ+Fp
uCPWQyBoJEiZqMdSDwrhmX8WSdS2r6TBT/K7QbG86o7GDN4yDBB/0frL/sUVL0UzQ9PycXgArpwB
wp1QPlNZbE60TJj4fovqB/ZLnfA60Mppg9GD8B9HU7/46auN0s263tBaTYH4eJDTx211FwXrPW1h
14aQETzTagHzKYBbyJvh9m7WQ54Uu5cb3i/ygEaJY/sH2nWMAIZ9ForBuHRccl/On5TWGF8rFSrP
QZqQ7nW4ttgcacnDJ0cekx+AiUgDJ8CE4ddY9NSuvQoj+eTtNk9PFS1tHB1RAHuYnilR5nG6U/Iz
6YLXh8GTLowz55Oevqo7cE+t8iR7C/WLOAUJm5I34Pn1FpK7rY0OaGWFlYKzeUKaplhp9Yqv+nwz
+vJjX8/5O1VY5sYyx/YjHNrwdKDvuvv6MXCt6oUQTrlT4JLdJZszndGN+nWsjL6irqbwoNxDAlr3
l3ta9fx3g3awR14JsYMBugSuP2k7d9pcLwYYcDq4SvPWN3F17xfI6Yj95oBZas1lG/poOqgzHr0D
c2gT9qKQtFSVqogusH5vYFAyf8tkKDgiausbR/Q7whj18KR0dRSeX/NLTR1rzafSxpa0mhRBQCN5
HYkN+3T1dSt2f0MQtliAe5xmHngnKV6myc5RotkiS8E/ruO+ve6kUqbKhvupOpaqa9go3kBeIH3B
m0U/2zWydsAxuhVpz9dAbOyLtKYEr5Zlt7OwyL6rPuUIIp/ai0d078kQ2zSlR8rxi/iHqjcRV9kC
dOikKkQDCyO1DA7vsDp0KTWYAiwSTj2F7GxOLO4+kRcQRn91AOs1HMg2/f0InTBOpwwmqPW+FODc
Bn4DKY/zt7suFcMyNTnqLBw8IOPXsGZmpG/hSr/mmTjsu/RiYVbhJsQ4OHQ+7OkXvJdKhs3XyQkb
YBFOzwM66I/QZ6BtobNAu+T2b03kFxWKfnJOBgStp5rh3ARnNgxNBdoPUKD2sgEpC9OmjfQ4osAi
w8O6R/ZXLV7tuCA/SOBLGXvJirPwq/VZHA/RmLwJ7L2C9XIeo/+W2DgaM981vgWYKPgl7ucoBuP5
HlK9WJca6DZ9H99/u78PKFQYdg5p9XCFL/ZYzT0jQCXDrTOkCXDL0iIfpSQZ99WUrE4sxXqIAci7
C9ra2Q4wh3eQU0EgClMWX6OYC8wfwYxqy3/NWNGA447w0x9q61Aep8qIbYasXJ0q+NrDYJ3TqL5Z
ngs66r1IH1bGtDeVe5hVfBoRkRg88/wyW+kr1FfCXdBRTYmgkPZY9sOrQvzr6BHKZaXI+PF9TJFl
sCfcT8yOern6hPydyMw5jRBgDaQF23gvtWn9Rjio+ITeQbePfTTuzKAL9RlLXfi1eUN7Yal2T8ph
K6eIphmEbKE/M0HeF7a+/PWx+Atqz3/iLNGgFAiuStKsydi5WIIsse/IUoGH+bdnycjqbKcZH/J6
HC8dOD+XptZ22p3vcqskTsY9syhq4HzCjOqqcveT1EmstgISkiYF/xVXx1xYROk2GeYv2w65ZV8H
7cHHZQ9zixUi5qK640RMI3PTsks/CLgBy2L43uDd9YQZyJWJs1duwSygcFrCjijU0z6BgUw+6IEr
LCbiS5NuGaRT76YT+HnW3gvBXlBXOAA1M7cIJxgYfhv/ih99XTSZXUJvIU3ArKpMFNAisj2uyR7Y
eWYHf3PE18TU/5X4H2l+zOoph72rLk+dCG5AGUyWSlkj4/jfmV2KAsXADbexGtxDxrCPEceJ7bF9
5gMpCkWzYru4AcN9a7SuOteNOcGmQ2n3HeUasvYdIXh0EmzIGj6iRRFGShR4c+AJnnhqjCsn7VEo
HXT4Bfn2dVd+8SGn0ADI8Lzex/g7wwIwrowTGesZSNuiWsiHIpDCFoe9q53nAt9fYpsF50J22Oym
KOcV46tgNJ99OzIs94LyAfiWPJW9bSi4Qu5iY+26m8/nFBbWJhgvAMQKSctHIJIxK3QrbR8FsSE1
46V0P2jX0CKXv6DS4wWJVTw2NdtVVyjF6XT4yvnkzcpBH5y2f7pI3Bcp567swx4djASfSpLVDh5m
JmHbvto6X+Zcb0jP5ofwGfKQi1MXy42Zo52l9rTYAZhLBOqqJfncFnGULKQ81VdAdfSO81+mL0Tk
U814BTvNjCWBgYvdmhlobrGuulhf6P8jUqUX6KLPiqLsKbcHk/dCVpYHg7tZ3sX1976DjA+tkufo
NI3Dt1wzMm0pcngkEYOhHvq/NksOvfsOoZp255CLm5/s9FWzO/bJsSOENs8kJEgqusPjBvztQs3C
jmVep7OXtLZ6wE9GCxKDPufNJrE+T98ko7xeckDCD77YfHsCUYWuacxh9XEuSepAz5F10PatCKcT
5jTNyT+ldJnxt9UGzUrquK101F2ZbhO52PQ8dHAKF0beVx/Ofj6T5lin7dwiRsmQW+AocWsgonEZ
paVS3cdCy0EdaOo+0/ViDbq16D1pm+gLnSWo4GPFD6/h5qwtsR+U/r1QrD+1hr3nFmAn2usQdrUH
DFME8i+uwY/7zLDNAMfx9YrPXZ2IwQ+PhbesuBr9ZcYFxrdNWyITJkDsySRpuWujT6T60Okr0iYI
mhuAUat7SmWbSQpy4qCJQYJ6Zir45CiinxkwgdsSR2w5dpTv+7SFmSa0h7r+SW4zq8qcI1OKufyK
jA3Oc0Kr//DLymZr4bTd+y3M68TiKIOZ2MPtlsJWQkcYklo97cY7g8wwVGguPGsiHsuqsAuAgEfp
Imxj4EBCwvvJKrUnljWHeqZgQQiflUCZWs1DaOCGIb2dyFUbVGIyBfVylx1XIzLYm3xQ+tZ62Inf
jG77wON30j7KkW47PKHxjuOcPDK7zNCiVvjLPGfxy2DcPXM4rEyD/fAcm9Qui+CYdRDrEiCU5QSq
k0nU6G/Jcag+j9ul8USRjON8S9HoPJwdMUL8VZZjRbbN66pqB2ze3UKhJD+iFxNOgbIFlp+ThGaZ
8HWp1SvinhtCL5nTbVAbxJqgusAUOdqXUmyadm8MmfCY1CT70UnM+/kBFvKl8RgWClr65jtl075n
srmPBSxAhW5JVSmAZ64fGBl8SZ0mWJataJxdNq2AI3WgGSOfZl56dkhgcD3/ngwF8oJ/jSF12GfN
JaVujrj00LhzYZNs3DNcm4QxDbRMzKW3wLkBPw6Y7W/As/UfNfWeztbi4FLSLET/7JFygNx7QKxP
x6k7q4zmcX7BNSIOlB5cqMC/jcLBzFuxSGnPxEOks/2KrKPnf7TD5XOTG6xfirdjDupkBy6t0q8s
c/lkE+Evc0lt4qSs6N2WLCaoqw9KB3fMEsaSIbHt9YbOlfkhFcQ6vjFXDCqf8VeGmRWkKrn6iccF
jxVXubFz9D2VOQoveVfTlTjRjiZOdf0o72oj/N7r/lOdFlp7HnNwG5Hv9hpEI92U2xsa8pCt8VPY
XeRpzY6LOksKhrLtba1mNEJMV44x5PfP1gvp98XofEAyYerMVvRqX0Ef4C4yCX3UvpWRkArSLvEn
3CsEtG512HT1fvqb3FPoBD+S91xfOQtl6yH+XXLVqxdp+2he/ifiJj4E3t19gvmqzWgUvKXhw2JS
Cj/iCOlRr6zl6vBS0Pe2UQ7DfrOWQ9gXrdJS36ISXCJ77DzKgKLPBF/GIJ80dU+zzTyB6CGN2WEs
FomkK3RwfTEy5wMsZRgfAke1JvmOEx+hftW1lBJ9I6h4yAX9aY50PqwSy4463n2CeSqPOWvZwcsu
IrzDRaLvza+YWo/QdS006p1dVY4HjtQ0QixoYHYdkQJdKusSv38BJfxqsDOYlxB6kODVQMBgaV/Q
+LyZd+ZNixMTkldfD50qNHhS+yZNQXVhZ26yMh/+aXfjDZ9bjAMJYIDNWpk37fjahyI3EVW6eCTD
asmyHZmx3wmJOZ36Ybzkg1gs8K2dDAyicA/eQbeVykPJiC6+k2aCDeZuuvyTOcVE42JfiZ7frsSk
57Kvkh37JyLhOx2g4SDLKlcsZCoCrWhjGNS3LuiRoJwGSnFwRZLx7dh6aq3lhMI4FcREEFMs/zN3
Os+K4oF8VMGnjLt69U9V5ulSSVIXKHMXCiyY45/ZIl4bYqdKI5zbU1hifmAIW93qIo+dEPUW1fMl
aSu7G4BRZkwhFWdau3tunUbILpUlNYfuZbtJkaAo5fTxRCVPhrbRS9gPoR0gGoVXQJi15+v3aThp
XQ+LyxaeRO06VXCQA7D57CLZhHB1ttlEoMlsj7+rWRinDB0648p3+VWOnDumvaJduXa8jwjd8+yf
KL/OufVM4kaa/z9H6k6cDa9LIh70nvjHYAyPPalycIPfuxJkybkuUwyq7nmM1nhzmCHI7MMj+ElA
Tf+PFUCK3UMVUBOR6x0QtN7PADMehPdloAVRxVymbVVZemMRFBBRxcGIcRRgfefjY6TJMVb2lef8
PYwwFxKU2a7eCMpfhx1jxcGT1hwIkuWTpHkR6K8eY++tU5N7Ms8VgSZ7nzWTSseqq6IBxyEonWux
u/WbhApsvZH3bkxEQ1whtJLT+YhuysJQbzWPvgK6AbCvxMET3j12xMhXqQgdZeQ/GGn7vPhLin2m
74FEXl4Sk2Oj0bj+UL6CVBp4czUqnjCjOOxs1/3E5L8P9Mgn4CVuAhelwsrL0uO8UIv7EfVIN20N
rIYU7F7DhTFsmxxmNWhI7CC/qnwDt0/qCuoVqe+arKocjgCldQULYPPgIjCLkw1+JkFI90v+bA6H
i6HGSOAwy+gw54uX08fj8iRB5yccsmXlEeDVHJpmzWjWzAtJCiPpjKX4pJ52KQch3Yw60rywQaZy
UnytgF+ch9W0xQ29sImZbjccYCmTNhB6zcsE2izEItBWGjy5PEg+W1YDuNSdGboXI6P72LCeOPWO
YODB5zRSiOeYp6XI8cqVDfMvB6OchJIIE0p9bI09OP9WpHGbC4yRRdASOP6WDkL7yQvEoXqmKPbM
0MBI86IXzqdenrLRLZPCXDRock6l7Jritk4M4I6VST3H/FS9PYlHaXEawfsYP/xTdc5PxfnLg3Ih
kjvao9XTBT1FjZ6joHjpzLZtpO9Ll/UKvcvw9kI3dQo+5qPpy+w+mKv4oTyvoWtj6/6Q9ll0llt/
V8RgNbjQ4uVSvp4wSIM9XadLU59/YK/r/pV3jy4xncznKszMWQNioUEi/4bYq7Wl/tD+tWjqA72C
bfp0jsgYbb1mDZ0HowJa9XjN1f9GdVWGMkCMEqDWkaokigU9YdAiP2yRk/TYU76NIkhbHFALiNi5
Je8oUzHyMu8szw5oGUcbF14D3Qwz76omSxoPWR0MdKirUR38keT2nI24QuGMDJ/MZwbOywEqOuqx
iR2D48VhttYEwnWz4bHimEu+ffRm+lyzhdGNeN1ZYTbmFj0JRot4xJYLeEAyte9aDdWnv29xLfKe
BN+MzR/GHFeXFCo85NLHk3XlaPA3OaRncWXmQo3F70NUQk5xl/JRd5z8H9ZJH4XOZ+2jcs/EIaZ3
npEKYnwWrx6BUJ8disCEaGgV1y1pj+5ipUKuu/quyZuGZqHXfa0Ul938nw7MhxSy72XHxRaJJX1z
Ek+FoMtHhjYp2nZoxTS+FiokVkFJnIsOVonv5FdZWTgNnDXVWcOr83wz2pHyR8vPnXgRM0l/BFWb
/2tOU9BMtltU6N2dNuXCjmYJq3HEpWhxBAKCObrX7XJZ9ebnmnc3BKHG0p6XrgHaG5iHwXncV7MO
0OsYpDLzrlhcAbqvK6D3dJHfL6SHPEqo0cG6KnUyiKoEy33e1cZ6Ri4do4x+w0GFG/Ao8xj5h67c
1UDcBx8aju9C3amNC3O2yxYKaoh9AVTpNNmMd4SYBlQ1HJCiUj3DE8Aroi91MJEYyNS8OK6mUkAd
S8w/cQFVPj4dcwAwijFMvt+yofR4Sz5X3g+6SKUr1ZU87qgaglu1h9EAOhdIttcV8WrTt4V/9RHh
VRqbGKeY2f4xJ1qTO4RDH7SNF4eZfI3BGAh+w4sQDp3MQnsfLf6p6ejTjjHoXCNEwTk3nurF2yVv
xtJic+HaDy3bCU3e44oHrDCElqZDrEKHOi7ofRKkzSgVuo1b0DbRY1MRhbdvCIiJlV1mpFJGldFG
LaLG4Y9s2FgrTz/RPM4CeRF674odR/9nis7w40C5hT9Tz+wvJo0Eim4E2+QhrZ2eDwYQYCeMeiR1
nhIjqs7qXih4QWzAlmR8gW390LG1MejqSzXq2He0Ye8Sf49gT68WP0Ukqr68hZD8bTJrjmIW3UJw
BH6u7gK+oU0tGXUevRpGJXeDjWs2B8U65GZq15tNaASPDazgqpyJ/b+hPx9XGynWLXYp+Wvj1AkG
l+kixskZGbznBABimjInTanEx++zIU6Ax+LV9ZHFXFVqgB8gWiRevB8FvPIYtHvVqfRvPZkgzuFH
TwwC/HcUImmfi4Poz4T8vY9h0Mxxxzjh87ggww4r8tTou5h/g6c6ACWb8WWEbTnJx/i/9js48LtF
tz7UmvVYAIGgXUYKwZyxJFOw4Oa5kTM9Fo5MayAlYjS35vfA/blCJknFVbYxECb6OytkdVQ/FU74
vIvm1GHqNFwb14lvopmO6xumUHqZUapP+1Qj9kXS49AtXYJq8gTsFfj2FhkmHY+6GNKciLyQNSi+
T1bMA6yJVsZUKr9FOblr3+pr8HeApDlWazbrAjW6EeAS86m+Gv2jk5yHRGqQPlloU+FaLVO4mx4X
gxditVbldL7Fn8B1HlwWt4Z/0jkiaGnlC+OgY3MVhtgzBGaamNP5jxTz03O6xECX3d38hmaa4Qrs
+yhoAT+EBtDVhwE0bB26fkGVIt0xlLStXKltuOA8q/mEDbvnP4MsE4n/CNVukAVcNNZOP0OvGQX7
Vfbm2zfEqg4zMeRluPPCeTKvaMLMFxLkfHl35wMMXJq2cd5crHjB/QtJR0lD/DRHlP2rEr2Gs4wo
ZQd+0k5eTks2lZNBrAAYSQFvEnVfjRRseTMc4LR5HnUR6m4I6BaprsD6bOHXFMuXVIQh6ofvHG+8
2Nppe+Odmz3xf6e65ZPkH7LsMz7FGv7mlTM/izf7/qjWCG4rxM7bIEnijuHWxQdyFk8NihtPmMzW
/dPDyyccoKBc72N9WC3TrWgUnUXALI6Rvqj8ZC8FV1+SzC5+w+IGjKcQXbXi4j9trN8s7kYJ8ijY
2bHyFrQ8k0pBIXXmXMmulzw9DGEsuisKzNplQN0qGsRnNtWAEkhe7s0/fLOLyWbQt2c9BlffHD/X
FFVPQIbU9UkSXbR0uwslTHaLt1jDZizCIZblouv169LN8KOF86rszp6w9UnPKcEulaGtA1TIW+6G
j6ujLqDU3zfPCFeNSv6Y+sgUi6pwhuwqsWHTbluvipHaUxDAqrYDE9h3ONeKB/AtKfyV+2Nitkyd
YXU4I9b+79WlseFmwaYbbKwCvzrY7iu8rsig1NnvsGHaJln+mNKaeahectWPk6OQ13aHLH5qdXaA
KurlizJMZZ5iihjrr37G/Yth6PynCtJDSO9z8xLdmJV+kqOillUY6UC527JnRvovGN9ZkaGJUbQZ
hlTP74pjmuwkq2UNenULnnuWpHbGU+t+775XeB9k6dB/fMGFModNaj1Bro0Q2/JyOXaW5y2XoFni
DFj/fUQrJIqT8+oju9aVoZE4a4PN4HAT5a3R1OdmVQoSnv/S+NNyyRCNPDVBabcsgfTKt/2x4F5Q
nSlXgr5/vSAgfdAL/CAch69voZ0d20SLBWs6M4bzx+QpO2URkfT+T3oBrkdmWwWOQmVM2ZE8nNmj
LHCcez3WJ4lO/HTtHBmxqTGQIrST9A4hyEO8uz41KSsk53WtrLhu7c/za78GL21+vPAPeRK7xwNC
1VGcNVmoMXlyFW6LCpUdI+4dNpaTdq9YaA1aNv3HZzWPe2qhUaERDlF+NlsShouByM2Cc3qXRVgK
uGn+9XqGJg3VmkLOxyp0BvKhcQNJ/RmJ8a8PvQLVAIm8M4jp/6ZwSRMCzeLAPvguy0VOjJiGiDez
DbUWJjQQhA+OyVK7F0Mih8NdU/A2JXtPEXs2aK5+EZ/0OuN1JTIVTKVyZT1jP4X8Jl4JhDiStCBW
ENq7nUZvzhWjjGSCAsI747Vfi6iD6xl4oB9hkz9+jpBpuMbCFDsliTCQy37IoWVgO9RSpy3UQyz4
lsS8sgt+ieIcXL5LZ1KWHGydkTGAH9vMBgBhVITuars9YlWjcckp+F4Y/D+NBvXoPjnh3Y1Eo07z
QjbrAHFHhmfRESdb0SC8Gn1ZZrhCT+GMMsMSkplSqNeUA/gD3o6FOn2Z74CrVs1es62j6TnYvK4Y
SXTTdq4HmkatKIjg0Yg9CVe1XAAq8wDVYWFlpFpV+61XhFPgP3zdl7XOni0cDmJ9/i2yD8QCzSAA
r+PANaabEe7mEyxC+V1qGYE1P8RglHBZeutRwLtQsld07E6/3mnRqUevDtUNeCU0XRkIkhJq4qDO
20jEIVrk9hXFZAacRCyv+NLbvBDkGwVMEmD1utY545Saraemxjy0u9tQHAnZWi1HDUHQX+2extC5
CDFHqRgDJhmJRMk5MGq6f/yR6czwyhTwzOTHdfnxeSCmZH2FZIc9tLq7f7bULSrmnThO8uBvXVwd
hbVzf03/qQziTavmhkNJPOy+paJq9a3So1ZmqoedFJk8telQjS7MHwaS+4dqD5sas6602n0PRsET
JHEljDQ1Rd+zk+ZZX/qUJsG2cU4rOU4y2H8WK3wA57RZKilO1POrnwxPpR750HwrJH2G17jlYF2I
pTteM4cygZhXprlUXlrytNWHGdVwgAHW/UQ7xhXMkdu6YBuX66H3p9HO3l8ao+ETzuBUa4yZZMB4
BXfO4VRV4b5fsvm/Jav1t+48Tw5GjCi949WUnABSVkMAosea08bcu1iiM/OXFcXuIATvKmpVTFRt
mI+NDFm9VjsZL5Nf89SVaq/XhlaIDvzRYucAj5jNUhl83yp0mqDanD7t+NpHJXZep8CKVQBThTA8
FSYr2Yu386Ly/dQOkKQo5w7R9H1xD0Rrv6LXCcDSuc85soT8pWHn9+Yl/kZncIiVirG+OhGnWhs+
qyLOMiFi4vgJGaJNuCmRkbhdIXDiBlleku924JJMpsRr9ugf2P8GTlDIS5q6S0upUOZbabU/n8ND
r3HoRYrJ87wW6qZ+lIZJQlS7EPRFlV3h2+8hBQbcpZcFuL1Ml4cu4l3NT29tIucG33E3xfs87gh8
K5O8ZD8q2kOJMtCoZ/BCorcaBwHuwMDLM2y6pRNqPpfnQwmu1lxzumcV0/Z1jYczhK7mbThZSg3B
b20AMduyguj8yCHni8UuKDERXFoBVnN4bDaE+4+AjUrlRVFcTRkpxmIo4KP4Ky/ShOx4j3Ssi6+v
/bXnzEZGVphGLjimLOTL+rRZe5wAyxN22H+L1ePLIIAu8bW1zCokAx0aKu9KvMi/Ruo+5lplyfsJ
ZAnfJBcXtJWHCImOPr9S/jJVA4MYeOOb0B9Wjlb3fk17CwD/vcveigv2heKmWQM3hNNYOJfZQu3t
lLwlElh68Jib6d+4fjf01tGtl/ZDJRjQq+OjzJAJyvuA7zRNeHXd+jnUYEgMPAjF/x3SPCCpe3RN
H5MU89kkqCSaNTAayIZ6hCs3N9Cq1txxV4M9PpJnGYRWUXQwHeJLmAzF0bw3/syxWwERBXOgx2gn
qG8Tf26iPvLGh/WryzOiGku4QEETUoqLTR7URgV6qSv62vhTV2mD6jgImklLYNUQFzPBx0KozjCB
hn/b2XLB8Eqs86YALmVV5PzFI3qIpUXul4SMVVIuXA9eQ+7g/51gASHfZ6YZQD154g+XGAKsN4OA
pZRfvN9KU5QKE/H+ek1n8VWjG4fH24dtg6BXfYr5Sef975ikvk0dHNvAfOrjhFh8kb6Z6kxkYwLu
I8LqUo3aLfsU5jU88o6oj+LVEi13blB/W79nqRI8RkurVeCtMZ0UYQsU6+m1IpyEd4Mupo4iT+z1
OO9aOfgH9cuNtaX72yFjrTDxBsoV36246T89vjA9EHx+ZhIPHt3F4tXjicWCU/lSsuBMYozo2zNe
Bl2jggU3hZheB59I63cvyf3u5oMjJlwBBl6Wd50xZwaXpfyaRb9t81514Z/mcg4FTrinTWT+aUkf
napdmZ/aj1qKw39nuXOEmcJKhRmrX/kS9YRrrvXZvUUJu1h3A9wRfzLAFdiu3hyRkaMiU2iKdkyG
A1j+1LODUKAJopaQ/GYgtpLUX0gHqmp7fVwueWPfsTBM0ItlFRDkc6AiJ+dDIpEd2zoQeE5qGShP
a8dFbk9aMHBYSZqmvND9tOAg4CAsKUeTldRrchewBOY1IL5joMlH11S3MRQzkBaSRXdZeDqIDDAQ
W/zZMUt+Gsvl9TiD4GCv4LOZyIRsNMHxavlneEiQ6GBw7wZ62khnPU/wTMY9qOxOmAyPKeVVz7j4
P39lW8pChrIOu0unQtB6mc6W5oFG1Bg5XoGpQslAAOo7tZkNinmEitlZU30oHiU/WR35AAwumBFA
EblQ3R3WT/sQQhpxcvtGZU79hRBe03BHQVRnEaOJeKSMmKlbKuXz11DzpW88gtSR+FbKXUYeSMH0
HhCv8Ie3AJNGoxNrFWo480yuZUUCBE5j+5+GZctTByxwhTA3EFheNORelIirhDnqYSYUzYBasnDZ
o/hcLCuRQj6Nf9CvebVNoUNVjh5ZFUBlv8xYgcyzvDVA9UlIu0vC6kSlHBwwxq45BZL+DtdiXmjh
zURsgvLEceWpB6Cha+6nuQli69O9gSQM/ttign//mYAXkjklxEsqoXA8UbCIT+IxKpZSO4KvOi5N
aCcqU/pofJmA0s4qXSD5uOK0MKeH7fcX3JRS1kCtxO973VDexOKXn2+maTioDS/ZAqtMcxqGAPES
72uuv44Fv5A2XWzolxHwVHv5BPbObXBZUPglMmWrYO6brJgVUR55O7HE6jxBcL/MmyBobFrvaHtA
kJWDaR6LzQmAyvsC4HhDNSWJ0HTaHWRS4UGfpM+kPZ1QT3EGeCZSg9ltH560P8YXHixTvummd7Gl
mfh6PVl3P+3PwVAGydhbndISUbxTDe92m+3MrTJALPKzf8A1nrCM77xIwPyHDtc/z+vth9fpZTK5
BwXhj1QGHSbxJbIKT2w8B5eOP9x8jj3OhD7dWjGLXLaXx5PeWtdu3xrZBJ4PMCtGjC2KOsNT3HRy
d7oKDprwxLscPz5c7Q6hoNghUzgpyLdgFVxTpN0H11jFO3s31sIcbye3RGW9FO/sKeDnwBjKlj1c
NoPm/Ep1VY7Sdarkfv8MUvcGkZfGsIWDkcUyzN4u4CJ7HqhRSHZpGwKvxG3G5/bnG4pruiI5wQC6
O3oiMN7l4b272CXJIRu4/1xljKMBdJECmEXMeUizBBGjvwgEglaHRZJlDqEcQW4dh2BDbbP4P79Y
Zc2NbMSPzPyC/ykfJrp9zLWzSvnyYO2CyeEBo3wei1LlSYAUVR3G87+ozoJBi9DKaixwZp84amXF
FaAW2isFG2NbEGm2Hx/A1aa/zP44S76NWaTlQoX+BNZXvQkX1ddiRy0y7Rugu2ipq5Zr11JSMPxn
9kjKDYrs73MGIQRJEwI3fk63XohwRSd1o8Jk+5NfCJS9L+KzAnfvW3OdmGFashyodLaCwc6q21CY
15IIAN9Z3yv4Y/yph6V1OHSpUHnhHSzVsozKk2uB4x+Jv/S1gj5oRFXfPxWkqdlfa5ZJwsYvaHXV
YLcqZIyQIQiVVgmb4RzvjtcJnd/7aPjNLM7LxjxnBvxtJzB91PntnfiKFcvFm/1XIVoKU1kxqXYc
1+/QyIb740NXKPIOfmKGEQxrpcRGXA3EHEbufF5v3aG8pZr01l27YzCcNPFQ0pHIEzC3B60zY1bG
yf2silb5fx3Vh8Z0C56oz77oKFqdFCtunAwIXm38wG3GvPluXxN5Vq9/ZtnMxAQkO49WzGsSX+s5
q83ljJGLOvIf/J5qunuz9SX17pqPVq8XP3k8TDNWIGTaWmU/xYXkGj53Q1u+vCnT804G37HpimgL
oykm9vSHSgIWlAwY/MJTRrCb/VNiQAGZwTZzJqH8AzntZhV5MkiNeWtLiTSdb2wyXrqB9TnNUhV+
dXVJMk1DpJ2+jnPbFaTx9hQztXFU7f0aJ4wuQQAKBDpJe5pr3wNEo6OZZZWSQM36AW0R5ffjIS+0
m0wbhtob+aqB7g4uXFNbVmr3E+Fsc3u50B6UPxCUmJriRUJ4mrmsuehe+AzEXWHKYruLB0/4Qh60
szmcJXfwko+07WNU5K+XhW10xbOiHamNBJ3D9r47ha2jjHvyOOIXhi3OUc+tT9a514lqCQ6v1yJ5
rtXTb/dxFxQ5toDUptbl3HHgDynW4IXHC68FmVWLK+20/ljUyxrIAXksSbAyw50JkcxBWPgpFybo
fyiaaAeZrO6VuXasqVNaY8LTdlXulOtGVCIVdXtdEUrmxN8AQmsSTCmvl3sh35eAoo5z04Q2ozG+
q3LfYDK7n72WdL8WsdGVdzRxlAF6pOyDUWKQu3BppMolvJWgB1jzJNuKoxbggyGtH6m4UD9zG/To
MduqVTE3Re/MQ1miyNb5YbOPFdvOLbN5LDesBvjc1zZitO3cNcsR+mkRbV3a/ZLga53Qud4mYhun
0pu43Df1n6QJf/YX5tYMxoG+obDFRLn52+ucS9odR/5kgPWBjj7/NvmDw/gq5fUvPolLQMbcitpI
6MqXIquBWTPUebY8UmdLMqaR2KRfe8IafgLphsJx1YOVgu50sorx/OxbLvcuBryNn5JYWLRF5vHG
Dhnn/hDLgiUp3CT0Bpj6IHYSwWm6OlYY89pmcNtAOqwJ1Rc2qAgXGI3WyfxIRMaOXtp6hiy6LLSa
i2BXWFm5X670OXrilRzFUHcytohvYZ4KEewflAvtCD/mf94iKXsLISVFsEaLqaqH7zFVl8m3KBHj
vEI3wNX6+nOlaj90Akwe3U5FJDfEuH5fpEUffgS3stFoz6C/NBnpsm2U8KPWaZIZ/Kj5zIswZa02
MaVvdVfUO710+OxcrBsZZB4ii1HvnlIGgdwfHMWIXmtKxj7X/mnHwn0OB7xCGe+TrwVi2EzUvR2z
tJS36e6wQb8JsprbzpPtOOyqUBa3K1AX0omtERLs8RD9Ldeib5dokOrkTy8BB7pL9/P/Y1ri7AIw
ICCVv6MZi28hPrIikQxXMiBUjYm5G8imKMCu2I/UMLiy9y5QZCxkwa4bvRCKaOfQ1d7CKtRWrs87
Ue8nCG+vs3Qo3HKffS4IZBnUHGsG++DMpNfSOZUxYRnpcf2Q3uPXCaRdB0GS4pXiFjyywsmb+POj
Pq2cZmuWAsOei8bOGh6ruSzkdc4UwkhfGIsVpHxm2wXItu8vJ+odiO3kHBDk1g0hqefcbQTIGXTY
+A2mxiBCwFRCja3eZOZ0fRxwV01CdNTR804y3Ta6+5IWQ2zIbRAkQffjhq3odjNW5uEE9IdLPvXp
2/Q1X6MsORmR4XsYVYeayiigxVXuAWs5gRs9oucFy4+P/mIVTVldzsp4iczwoYFVlSzPUmR4Awj0
+rjV8zaB7sYvpiid8SgG9XWh+LqXi2qv9BPzb1Y1fLAODQr8rmx6/MeZfMqrLtKnhtjImW5PxwmW
JTr4d1Ymmrr16m9DutzuMbFLOJFMslnDdGd6uywmy8VedwXMKZo2m4JbPmNqXPVMP/8grXiarXqs
Vcr5H1ltW275Swo30YK7RUSlYCqLQIsKLXXferDmZcWgL9FXhWT/H/M02MvwdAyKEvcQkTwRNIXf
2kefbq5u5JoPx9SDTIXmw5EseAqv489eOdwsV8vkhXQQfpU/oOAMEOiu85l9TpMl3rfl1QmSTIwS
X6J0C8puMiz5AnsLLQvWJZUb5JZ0u+iinsx74upsuetFpNura14k2gDB6XcaFY3Gu0e051YVbBSF
3nF/4LxbGIcCVxaGmrld51Pr3wPKgvWNXOMiBSijijfJ3ZQRUfNTf8IGpIVX/Irfq8bAuH2RHm/S
6ZtPR/PE8/Ly10W4G/1WfX4tTK0PrfGaddIQlgFSMjnk9rT9phZG8qvUO+OeBi3R69tQVY+Ujw5r
5aSlMgOyRVDB4uRHas3QaxJu1iY/iNafLMyPObPnfrEhW3zfiGxC+DDz9y9Npx/pevrkou6cpHZD
YsSNuMgd+l0iHmlWG12WkC6xQaiqQx7pN2t7XQK81E6z0I2UubB5/FaobHVy8F9EQc7kaUvU7jiJ
O2ewtQvW5L/HncMZnfpdH1Zgu/9w/bLkXOUppnCCACtROzmOuHqh+FVGY7A0U6eClKqbmNhuu3kE
AR4VBbgd+IrCNVwilqWG8k+05qvHYB70Fn26Usl9L/hHcJejMfZpZ2D2A9S7IypUli92ZPcNRpdp
lkSE1hRXnLo0BeOITXaP/jLSgxn9ngjzQljO0AAhTcE+xUJgC7dsBMh7kUjFXsVVUSIAxBeIau7Z
fjpr4tSToEBUcfLzx/vkKvcpdxxvmWwqBm9zEoA8XDkDPWLfk9IttkmYni8x/z2QetU3qdqN790t
Udtywl4oGZrQiiMD6d9SBiksbLhUQjpgpcwug0SFRRKP6qiAfX26jQjIJsHWh9HtET6uWTf16PFv
qbAIPSJiOE4Ds8wQFRRw06N9blvimhgEX4DvYZ8jr1Ktitf3mhp7KyQa2YcwKGmzchNA+YXEqah4
1UhwJtRdst3xKmH97bcQ2gnk7/jZ4s5n+yAP3kBoX5Yzmx4S6+fsg966lRWcdKhcfL8oggPakeM8
Ezm81ORFdX39W3k6JPVFsW10ZiILpevbKsIx2xRSIsmWqnbSPIa85UkjDJvGkNXc+HqugjEsGjkj
matd85xHcCbCAkWFmpM/CD6g6XXLjjgxeMyjVa5QkYQDXbMAyIGPaqABsJPzRM23guhZU8DfIZjl
wNRIEL12V+mGgpT6a4yFobwpvL6Fjv/Otlc2WKb83CW7kCjHGlEXgUvbWVxFTUZetPE8y1SPPXOq
sRznJC/W9D9ePHBhy950kyt2R9BA6NasghoYAEv+edFpbM/MfvInVLSOQ2SBwiFCV4FL0FToQjHB
PffZ/PDuIGMXbyG1YBk1jhQQGqkk8SO7hZXL2bplV6/M0MIKow1ucn7Uqn/pFaYLxI5XAG83e5d8
BPSh4gOEbtfqj3AtvJI0TkajjAzDmYMlWiZj2hNbwRTZvRH2XzsGECoCWncX49oADQ/sGAbF5N2H
sW5f+zGa1DD/HxvG8RKLA/dl+1SiWxv2xOT6Fp94nqGVL0508W5H2+Eb5Db9x+mWkuPZ35zzfn2X
oPgj1vq5nEdvxlCyvsgyaoKCo4cjK5ry8055HnB717gKRed1XFaj1BVYWctKUiIOL7OsDpYDn7UD
rbylZyPF53zXtN3S1o6BploNz1bqjzhkCW53PPVTWjFh5htVVFlBb7xN00mdJ7Vo0IYNz2yIRA33
C8VZoGxw+SguwHh0+UPsqtEFjVit2SW5mFF3u+9bKUJ43CaySmZjJUc6pHbEOMXksmaWn/QYjktb
XH/xoRT/vDXcoi0NYJucy8ojX8DRB/60pW38WP23IPvHTH5KLXRGI1VCvfhfg6gLwTz3mct7JAT5
DfJd46SmoMWhhCBVeEE45cuBV+wW5gaVYfBwIjRGrrgCSf3lwRvwJEKNZtzFkrOJi6PTE/958nvc
nm0taHNtHNXm0dLq/NaO9fmxZVjaocFTJBwgI7wSeZfIbzZz4VrtmCtLzzXKcOcfSAtXPh7Di3ce
CgbvcN6bB6wuakjeoe7j66zrO97B8GLbYltARu4eMmZOgLvVogau9UKVewhUqg6u12WfpfBwjCnX
ULqMulNta/+AmkP2LskaLfyDX0C+rPG58Dq8DCtFjaFlLGKHDtVeVjYfo46bP4vbbgxCTAokIni1
9gjvW/6hyrObOfV1ie+qmZitij96zzDhE3KTYlDipjtPkDdDxMzXQENLiFicBDQTAJqASo7MjSDh
LSFY+pypFOLOlznXAJ60UMelx8bhBTia3mkLrzxuV3l6E2JlktHWJ06xoBeViKekLbugIozxJ4tA
O3lCZphAPRyet+1RdACCIKkObnBwJAsilvSiTJpqCBtjw+hUBAkpYPasOzYiNPfTb65nUqU0bNJH
9JSPYUZ1Ha/w27qdGsQ19zJhXvHfMV5m4K6qVzSNhaanmpxd2MsH2QFLhBMfIvfZqbbnhmpKdyVo
/IGXQgwikic67UxqOFaiZ832S+uh9Vva2sKhE3FswzpHi30Busl+902uzsSKKZ2D6kO1FBGs+I13
v33M6TFnyOFL7FTu1/pCSYAooWfouCVfN/KamghT4ur7iV4OurdoeWa2XFLYg8Z0iF3D4r2WlxU9
rhimSjMIdV6HyITtTWiVWXwD4w1n4KFf3UlxlgJuqCmZ81P0Z5qP2oCFYAd+dhNSJbF0T30JZTVN
gIOrnS6lhbJt7y30ITIwlo4bwps1gTQFyOvlZOuXouinl0t2fsK/k0vcuCMNHh+TP21HteJYWRxv
pSuTF0K1rISeeHcvkVt/L1oa3s45bQJDXLOSy4RbydMbofj9NkBU0Tf0/TQ/G+M4Q9jGUhnWRcSH
PZ5FD5b+6/4WzifJa9v2PlvFIAvK4GDEr5seKRz+99qdPYXSYTPDrByN8xjO9h0qy9QUa9k2x8ik
D2yLEuHxm/2/oDrP1znB/XzXs+wqsR9nPt83++/1BcTVo+1GZ0hgdvheQFVJrK1+Oz3vX6wrjjhd
z9AuBk3EmJOiPGuaSAsWIy65c53IHNOTPiN5qyY725YsFhggLPRoMnmEYLhrF7hzmrHJIli32338
5VPJzspKLVKh6zt9UwNA6GlwsU3T4sjhyKiz6SqW56Adkg7AKTpWy5Egz1zEHrLTgJIreW+ljgOm
1Z9sPDx3ignHe+d2bWMxj9YwWDA/2QFIxskGU3UO0iyZrrnN0FghiInbX+qDcJ6oyR/ZhXmN6Ut2
BHQjLKLRU6oID1/JsT5O17AgkplQ2kRcdr8/ZT9W07TUsn5xy2To30rt7yeZ4gAktqGt0k3Oc0TK
L/AtryxpyhriOoaKDQYwubvACkrGoijU+L8uM/er2RIicSdWI6ITmBQGatrT6ZtFtB4486HOREBR
lQF9EWykfYHwhm2iCq8uyaCVHwfIotTj4EqvQRQo0HVoa0pP+mEN5IZWJgyJ00f/GVz3UyKLrKby
XwMyESiY+fCDtDA/c2swg6pXqPArMSDkgyXx1m7RuBrfUNbKZSSpnaYhlroh2mWa1BQom6gKy2pI
skU+pKxX0jhZFvFpcZ9QbIWfNqeqE3qgEjf0EKFrdbrL+8J/Oqsd6NmAZPMhgZl1ygUrzgAq8CrK
nFazLvhvVt98nNg68Yx6WVHXUucfK3nSc8ytIz8c/dPlI14VcjCHHSZ0mX+8eW5A61U28V4xPJ9g
D8NbOc/ZzURJ7XMstvYMzXtfC51N0nTeiXpTn8lVe/LNZ2JDhnem3SUnU+gfKTwHUquD1XKF/1AB
jyN7xUwO9QwT854ATgTWGLoVBvnzf09+iK/OPU5RzMTOiHeJ1fgWc0V3JceyuOjS252oJKip9vB8
qYJoVmWsneuwIhmKXVjnredmOoj5kya1OsYwkRqwRHm7O+teJ9XxMr9cx/nByxLjp3XP6TnuO8Tx
tQ7Cz/R6RS0a0em4e9EBV4VY4B6aSMzWg1chotYC/Rjv3vcT1exQdaJWXEZbpyDgjg/rwQ+r4c2k
tqmgIC4EK9evAZobD75O4vkJGC9HypjO0Kwsa72Am52sXjPArA27ckh304vPfq9AquRKW1RbR/KG
Ysjv4vRTfWIqoMJbVZ+D0NG+U1xPH40U/NG5+Q7mFh2OLNv7UDe/V9h4N2181ZWAEOmzv4zxQvx2
Fvn5sF2aJsPZ3eIBOc57RcmXbVWcnR6yB3ZWqYLAB+xKufc34S+tG/Y1nIjIKTNGzBYYZOD5RHiK
gDD84g/8L5w7OVL3p9LJBeKK44faXI1x6/aOcaBuc3iKfFOE9C2f3vmMdRhGAg3pOEgoBs+V7ykE
3XO97QpJ74meo2zaj84nqy/iTWdK1+YnaC19LVC1nITkHJhLsnU1INacyUdKRCGpMEXyhus1hRUV
uwIInUavtLQzt4bjLN03wLIWcNIHGr6DOIFBq8rQXx4Ul0UoAkYfH7RsvHbKR+0CXbgrWwSrJM5A
vJgRDgmXl1gi4Lcs2xoXwktJccmJwonKck6roeQOhml0Gcrgxue+zERuJyi3LGUKd5CISS7ZqSPc
4xjXfc+MmuBHpavpiI/2Ax7cNNhWllRo179c3uDRAPQQx2esHlXe4TDATMkwILCfAgbQpzLbgzGH
fvuzLv3YeiB1Zt4FrHjuaUgO2X3hoEBNLzK23QUYGQts1QPuN6Gc26V7ZEKoU9cWqF66Z9jglHIp
Ns7yPUw8Qgfhbu/FmNh++/v3bZQGsN8X2HB98LIUL+5PV8SdiFZgrD0S8am55+5VUV/dc2gctfjA
XtJ2n6tSdcPyaCQ6pLLAhjgUM7eDd0q4vd3DNBrAxAsHvD2q4J92XBSek1BkjkxaBtkoGuFIefmP
ygUKVW0anlRbYSm+ctoVRDnmkJjNpQ23ZRbeZXeVuneJGwxQlXkaSMoYcP6gulzxhYsV4HI6+CF8
NQAaDYb0UaliMRG3HA1byXnPpIuMd8rDcydGi6QNidwR49uEIpI8ooxRYLiRGIvbkNo9fUtr7hZb
Ws4N34eTs/HOi8TJsQ28xSGEwjqd5EfnXQ==
`protect end_protected
